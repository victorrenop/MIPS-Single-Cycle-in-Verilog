
module BIOS #(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=400)
( address, instOut, clock, autoclock, rst/*, changeSource*/);

		//output changeSource;
		input [(DATA_WIDTH-1):0] address;
		input clock, autoclock,rst;
		output reg [(DATA_WIDTH-1):0] instOut;
		reg [(DATA_WIDTH-1):0] mem [ADDR_WIDTH-1:0];
		
		initial
		begin : INIT
			mem[0] = 32'b00000000000000000000000000000000;
			mem[1] = 32'b00111000000000000000000000000010;
			mem[2] = 32'b00110000000000010000000000000000;
			mem[3] = 32'b10011000001000000000000000000000;
			mem[4] = 32'b01111100000000010000000000000000;
			mem[5] = 32'b00110100000000010000000000000000;
			mem[6] = 32'b10000000000000000000000000000000;
			mem[7] = 32'b00101100000000010000000000000000;
			mem[8] = 32'b00001100001001000000000000000000;
			mem[9] = 32'b00110000000000010000000000000011;
			mem[10] = 32'b00001100001000100000000000000000;
			mem[11] = 32'b00001100100000110000000000000000;
			mem[12] = 32'b00011000011000100000100000000000;
			mem[13] = 32'b00110100000000010000000000000000;
			mem[14] = 32'b10000000000000000000000000000000;
			mem[15] = 32'b00110000000000010000000000000000;
			mem[16] = 32'b00110100000000010000000000000000;
			mem[17] = 32'b00101100000000010000000000000000;
			mem[18] = 32'b00001100001001000000000000000000;
			mem[19] = 32'b00110000000000010000011101011000;
			mem[20] = 32'b00001100001000100000000000000000;
			mem[21] = 32'b00001100100000110000000000000000;
			mem[22] = 32'b01110000011000100000000000100111;
			mem[23] = 32'b00110000000000010000000000000000;
			mem[24] = 32'b00001100001000100000000000000000;
			mem[25] = 32'b00101100000000010000000000000000;
			mem[26] = 32'b00001100001000110000000000000000;
			mem[27] = 32'b00110000000000010000000000000000;
			mem[28] = 32'b10010100000000010000000000000000;
			mem[29] = 32'b10001000011000100000000000000000;
			mem[30] = 32'b10010100000000000000000000000000;
			mem[31] = 32'b00101100000000010000000000000000;
			mem[32] = 32'b00001100001001000000000000000000;
			mem[33] = 32'b00110000000000010000000000000001;
			mem[34] = 32'b00001100001000100000000000000000;
			mem[35] = 32'b00001100100000110000000000000000;
			mem[36] = 32'b00001000011000100000100000000000;
			mem[37] = 32'b00110100000000010000000000000000;
			mem[38] = 32'b00111000000000000000000000010001;
			mem[39] = 32'b10000000000000000000000000000000;
			mem[40] = 32'b10010000000000000000000000000000;

		end 
		always @( posedge autoclock )
		begin
			instOut <= mem[address];
		end
	
endmodule 
