module ControladorHumano (OPcode, hdt, RW, MW, RDst, ASrc, MTG, PSrc, Jmp, Jr, ALUop, halt, flag, out, MO, Jal, hdFlag, writeInstruction, setProcess, menuWrite, changeSource, changePC, changeContext, bw, BSrc, tw, tr, tb, rwc, MWC, uart_flag, uart_write);

	input [5:0] OPcode;
	input flag, hdt, uart_flag;
	output reg RW, MW, RDst, PSrc, Jmp, Jr, halt, out, Jal, hdFlag, writeInstruction, menuWrite, changeSource, changePC, changeContext, bw, tw, tr, tb, rwc, uart_write;
	output reg [1:0] ASrc, MTG, setProcess, BSrc, MWC, MO;
	output reg [4:0] ALUop;
	
	always @(*)
		begin
			case (OPcode)
					6'b000000: // nop
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'bxxxxx;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							changeSource = 1'b0;
							setProcess = 2'b00;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0;
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
 						end 
					6'b000001: // halt
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'bxxxxx;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							halt = 1'b1;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
 						end 
					6'b000010: // add
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							changeSource = 1'b0;
							setProcess = 2'b00;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
 						end
					6'b000011: // addi
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							changeSource = 1'b0;
							setProcess = 2'b00;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
 						end
					6'b000100: // sub
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00001;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							changeSource = 1'b0;
							setProcess = 2'b00;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
 						end
					6'b000101: // subi
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00001;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							changeSource = 1'b0;
							setProcess = 2'b00;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
 						end
					6'b000110: // mult
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00010;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							changeSource = 1'b0;
							setProcess = 2'b00;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
 						end
					6'b000111: // div
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00011;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
 						end
					6'b001000: // slt
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01010;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b001001: // shr
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 1'bx;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01001;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b001010: // shl
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 1'bx;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b001011: // lw
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b01;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b001100: // li
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b001101: // sw
						begin
							RW = 1'b0;
							MW = 1'b1;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'bxx;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b001110: // jump
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'bxx;
							PSrc = 1'b0;
							Jmp = 1'b1;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'bxxxxx;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b001111: // jump register
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b1;
                     Jal = 1'b0;
							ALUop = 5'bxxxxx;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b010000: // xor
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00111;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b010001: // and
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00101;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b010010: // or
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00110;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0; 
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b010011: // not
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00100;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b010100: // xori
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00111;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b010101: // andi
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00101;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b010110: // ori
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00110;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b010111: // beq
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b1;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01100;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b011000: // bneq
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b1;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01111;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b011001: // beqz
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b1;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01100;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b011010: // bneqz
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b1;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01111;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b011011: // bgt
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b1;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01011;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b011100: // blt
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b1;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01010;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b011101: // bgtz
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b1;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01011;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b011110: // bltz
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b1;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b01010;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b011111: // in
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b01;
							writeInstruction = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
 							if (flag)
								halt = 1'b1;
							else
								halt = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b100000: //out
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b01;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b1;
							MO = 2'b00;	
							writeInstruction = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
 							if (flag)
								halt = 1'b1;
							else
								halt = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
                6'b100001: //jal
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b1;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;	
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b100010: //cpyHDToInstr
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b1;
							hdFlag = 1'b0;	
							halt = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;				
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b100011: //srprc
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b01;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b100100: //src
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b1;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b100101: //swprc
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b10;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b100110: //smenu
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b1;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b100111: //memhd
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b1;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
					6'b101000: //loadpc
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b10;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
						6'b101001: //changepc
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b1;
							changeContext = 1'b0;
							bw = 1'b0;
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
						6'b101010: //lint
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b01;
							MTG = 2'b10;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
						6'b101011: //ctx
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b10;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b1;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
						6'b101100: //ltb
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b11;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
						6'b101101: //stb
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'bxx;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b1;
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b1;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
						6'b101110: //hdmem
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'bxx;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b1;
							BSrc = 2'b01;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
						6'b101111: //stm
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b1;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b1;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
						6'b110000: //rtm
						begin
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b1;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
						6'b110001: // lwc
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b01;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b1;
							MWC = 2'b01;
							uart_write = 1'b0;
						end
						6'b110010: // swc
						begin
							RW = 1'b0;
							MW = 1'b1;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'bxx;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b01;
							uart_write = 1'b0;
						end
						
					6'b110011: // send
						begin

							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b01;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							writeInstruction = 1'b0;
							halt = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
 							changeSource = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b1;
						end	
						
					6'b110100: // recv
						begin
							RW = 1'b1;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b01;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
                     Jal = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b10;
							writeInstruction = 1'b0;
							hdFlag = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
 							if (uart_flag)
								halt = 1'b1;
							else
								halt = 1'b0;
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0; 
							BSrc = 2'b00;
							tw = 1'b0;
							tr = 1'b0;
							tb = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
							uart_write = 1'b0;
						end
						
					default: 
						begin 
							RW = 1'b0;
							MW = 1'b0;
							RDst = 1'b0;
							ASrc = 2'b00;
							MTG = 2'b00;
							PSrc = 1'b0;
							Jmp = 1'b0;
							Jr = 1'b0;
							ALUop = 5'b00000;
							out = 1'b0;
							MO = 2'b00;
							Jal = 1'b0;
							writeInstruction = 1'b1;
							hdFlag = 1'b0;	
							halt = 1'b0;
							setProcess = 2'b00;
							changeSource = 1'b0;
							
							menuWrite = 1'b0;
							changePC = 1'b0;
							changeContext = 1'b0;
							bw = 1'b0;
							BSrc = 2'b00;
							tb = 1'b0;
							tr = 1'b0;
							tw = 1'b0;
							rwc = 1'b0;
							MWC = 2'b10;
						end
				endcase
			end
endmodule			