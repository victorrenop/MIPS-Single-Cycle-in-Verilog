module InstructionMemory (adress, InstructionOut, clock, autoclock);

	input [9:0] adress;
	input clock, autoclock;
	output reg [31:0] InstructionOut;
	reg [31:0] mem [180:0];
	integer flag = 0;
	
	always @ (posedge clock)
		begin
			if (flag == 0)
			begin
				mem[0] = 32'b00000000000000000000000000000000;
				mem[1] = 32'b00111000000000000000000000110101;
				mem[2] = 32'b10000000000000000000000000000000;
				mem[3] = 32'b10000000000000000000000000000001;
				mem[4] = 32'b00101100000000010000000000000001;
				mem[5] = 32'b00001100001001000000000000000000;
				mem[6] = 32'b00110000000000010000000000000000;
				mem[7] = 32'b00001100001000100000000000000000;
				mem[8] = 32'b00001100100000110000000000000000;
				mem[9] = 32'b01011100011000100000000000001110;
				mem[10] = 32'b00101100000000010000000000000000;
				mem[11] = 32'b00001100001111010000000000000000;
				mem[12] = 32'b00111111111000000000000000000000;
				mem[13] = 32'b00111000000000000000000000110100;
				mem[14] = 32'b00001111110111101111111111111101;
				mem[15] = 32'b00110111110111110000000000000010;
				mem[16] = 32'b00101100000000010000000000000000;
				mem[17] = 32'b00110111110000010000000000000001;
				mem[18] = 32'b00101100000000010000000000000001;
				mem[19] = 32'b00110111110000010000000000000000;
				mem[20] = 32'b00101100000000010000000000000001;
				mem[21] = 32'b00110100000000010000000000100111;
				mem[22] = 32'b00101100000000010000000000000000;
				mem[23] = 32'b00001100001001000000000000000000;
				mem[24] = 32'b00101100000000010000000000000000;
				mem[25] = 32'b00001100001001010000000000000000;
				mem[26] = 32'b00101100000000010000000000000001;
				mem[27] = 32'b00001100001000100000000000000000;
				mem[28] = 32'b00001100101000110000000000000000;
				mem[29] = 32'b00011100011000100000100000000000;
				mem[30] = 32'b00001100001001010000000000000000;
				mem[31] = 32'b00101100000000010000000000000001;
				mem[32] = 32'b00001100001000100000000000000000;
				mem[33] = 32'b00001100101000110000000000000000;
				mem[34] = 32'b00011000011000100000100000000000;
				mem[35] = 32'b00001100001000100000000000000000;
				mem[36] = 32'b00001100100000110000000000000000;
				mem[37] = 32'b00010000011000100000100000000000;
				mem[38] = 32'b00110100000000010000000000100110;
				mem[39] = 32'b00101100000000010000000000100110;
				mem[40] = 32'b00110100000000010000000000000001;
				mem[41] = 32'b00101100000000010000000000100111;
				mem[42] = 32'b00110100000000010000000000000000;
				mem[43] = 32'b10000100000000000000000000000010;
				mem[44] = 32'b00101111110000010000000000000001;
				mem[45] = 32'b00110100000000010000000000000000;
				mem[46] = 32'b00101111110000010000000000000000;
				mem[47] = 32'b00110100000000010000000000000001;
				mem[48] = 32'b00101111110111110000000000000010;
				mem[49] = 32'b00001111110111100000000000000011;
				mem[50] = 32'b00001111101000010000000000000000;
				mem[51] = 32'b00001100001111010000000000000000;
				mem[52] = 32'b00111111111000000000000000000000;
				mem[53] = 32'b01111100000000010000000000000000;
				mem[54] = 32'b00110100000000010000000000000010;
				mem[55] = 32'b01111100000000010000000000000000;
				mem[56] = 32'b00110100000000010000000000000011;
				mem[57] = 32'b00101100000000010000000000000010;
				mem[58] = 32'b00110100000000010000000000000000;
				mem[59] = 32'b00101100000000010000000000000011;
				mem[60] = 32'b00110100000000010000000000000001;
				mem[61] = 32'b10000100000000000000000000000010;
				mem[62] = 32'b00001111101000010000000000000000;
				mem[63] = 32'b00110100000000010000000000000100;
				mem[64] = 32'b10000000000000000000000000000100;
				mem[65] = 32'b00000100000000000000000000000000;
				flag <= 1;
			end
		end
	always @( posedge autoclock )
		begin
			InstructionOut = mem[adress];
		end
endmodule
	
