
module HardDisk #(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=4400, TRACKS=2)
( clock, autoClock, track, trackPos, writeData, readData, hdFlag, rst);

	input clock, autoClock, hdFlag, rst;
	input[(DATA_WIDTH-1):0] writeData, track, trackPos;
	output reg [(DATA_WIDTH-1):0] readData;
	reg[(DATA_WIDTH-1):0] disk [(ADDR_WIDTH-1):0];
	
	initial begin 
	/*disk[0] = 32'b00000000000000000000000000000000;
	disk[1] = 32'b00111000000000000000000000000010;
	disk[2] = 32'b00110000000000010000001101010110;
	disk[3] = 32'b00110100000000010000000100101010;
	disk[4] = 32'b10000000000000000000000100101010;
	disk[5] = 32'b00000100000000000000000000000000;*/

			// SO
	disk[0] = 32'b00000000000000000000000000000000;
	disk[1] = 32'b00111000000000000000010100110010;
	disk[2] = 32'b00110000000000010000000000000000;
	disk[3] = 32'b00001100001001000000000000000000;
	disk[4] = 32'b00110000000000010000000000000000;
	disk[5] = 32'b00110100100000010000000000000100;
	disk[6] = 32'b00110000000000010000000000000000;
	disk[7] = 32'b00001100001001000000000000000000;
	disk[8] = 32'b00110000000000010000000000000000;
	disk[9] = 32'b00110100100000010000000000100111;
	disk[10] = 32'b00110000000000010000000000000000;
	disk[11] = 32'b00001100001001000000000000000000;
	disk[12] = 32'b00110000000000010000011101010111;
	disk[13] = 32'b00110100100000010000000001001010;
	disk[14] = 32'b00110000000000010000000000000000;
	disk[15] = 32'b00001100001001000000000000000000;
	disk[16] = 32'b00110000000000010000000000000000;
	disk[17] = 32'b00110100100000010000000001101101;
	disk[18] = 32'b00110000000000010000000000000000;
	disk[19] = 32'b00001100001001000000000000000000;
	disk[20] = 32'b00110000000000010000000000000001;
	disk[21] = 32'b00110100100000010000000010010000;
	disk[22] = 32'b00110000000000010000000000000000;
	disk[23] = 32'b00001100001001000000000000000000;
	disk[24] = 32'b00110000000000010000011101011000;
	disk[25] = 32'b00110100100000010000000010110011;
	disk[26] = 32'b00110000000000010000000000000001;
	disk[27] = 32'b00110100000000010000000011010110;
	disk[28] = 32'b00110000000000010000000000000001;
	disk[29] = 32'b00110100000000010000000011010111;
	disk[30] = 32'b00110000000000010000000000000001;
	disk[31] = 32'b00110100000000010000000100001101;
	disk[32] = 32'b00110000000000010000011101011000;
	disk[33] = 32'b00110100000000010000000100001110;
	disk[34] = 32'b00110000000000010000000000100000;
	disk[35] = 32'b00110100000000010000000100001111;
	disk[36] = 32'b00101100000000010000000011010110;
	disk[37] = 32'b00110100000000010000000011011000;
	disk[38] = 32'b00101100000000010000000011010110;
	disk[39] = 32'b00001100001001000000000000000000;
	disk[40] = 32'b00110000000000010000000000000001;
	disk[41] = 32'b00110100100000010000000000000100;
	disk[42] = 32'b00101100000000010000000011010110;
	disk[43] = 32'b00001100001001000000000000000000;
	disk[44] = 32'b00110000000000010000000000000000;
	disk[45] = 32'b00110100100000010000000000100111;
	disk[46] = 32'b00101100000000010000000011010110;
	disk[47] = 32'b00001100001001000000000000000000;
	disk[48] = 32'b00110000000000010000000001000110;
	disk[49] = 32'b00110100100000010000000001001010;
	disk[50] = 32'b00101100000000010000000011010110;
	disk[51] = 32'b00001100001001000000000000000000;
	disk[52] = 32'b00110000000000010000000000110010;
	disk[53] = 32'b00110100100000010000000001101101;
	disk[54] = 32'b00101100000000010000000011010110;
	disk[55] = 32'b00001100001001000000000000000000;
	disk[56] = 32'b00110000000000010000000000000001;
	disk[57] = 32'b00110100100000010000000010010000;
	disk[58] = 32'b00101100000000010000000011010110;
	disk[59] = 32'b00001100001001000000000000000000;
	disk[60] = 32'b00110000000000010000000001000111;
	disk[61] = 32'b00110100100000010000000010110011;
	disk[62] = 32'b00101100000000010000000011010110;
	disk[63] = 32'b00001100001001000000000000000000;
	disk[64] = 32'b00110000000000010000000000000001;
	disk[65] = 32'b00001100001000100000000000000000;
	disk[66] = 32'b00001100100000110000000000000000;
	disk[67] = 32'b00001000011000100000100000000000;
	disk[68] = 32'b00110100000000010000000011010110;
	disk[69] = 32'b00101100000000010000000011010110;
	disk[70] = 32'b00001100001001000000000000000000;
	disk[71] = 32'b00110000000000010000000000000001;
	disk[72] = 32'b00110100100000010000000000000100;
	disk[73] = 32'b00101100000000010000000011010110;
	disk[74] = 32'b00001100001001000000000000000000;
	disk[75] = 32'b00110000000000010000000001000111;
	disk[76] = 32'b00110100100000010000000000100111;
	disk[77] = 32'b00101100000000010000000011010110;
	disk[78] = 32'b00001100001001000000000000000000;
	disk[79] = 32'b00110000000000010000000010000111;
	disk[80] = 32'b00110100100000010000000001001010;
	disk[81] = 32'b00101100000000010000000011010110;
	disk[82] = 32'b00001100001001000000000000000000;
	disk[83] = 32'b00110000000000010000000000110011;
	disk[84] = 32'b00110100100000010000000001101101;
	disk[85] = 32'b00101100000000010000000011010110;
	disk[86] = 32'b00001100001001000000000000000000;
	disk[87] = 32'b00110000000000010000000000000001;
	disk[88] = 32'b00110100100000010000000010010000;
	disk[89] = 32'b00101100000000010000000011010110;
	disk[90] = 32'b00001100001001000000000000000000;
	disk[91] = 32'b00110000000000010000000001000001;
	disk[92] = 32'b00110100100000010000000010110011;
	disk[93] = 32'b00101100000000010000000011010110;
	disk[94] = 32'b00001100001001000000000000000000;
	disk[95] = 32'b00110000000000010000000000000001;
	disk[96] = 32'b00001100001000100000000000000000;
	disk[97] = 32'b00001100100000110000000000000000;
	disk[98] = 32'b00001000011000100000100000000000;
	disk[99] = 32'b00110100000000010000000011010110;
	disk[100] = 32'b00101100000000010000000011010110;
	disk[101] = 32'b00001100001001000000000000000000;
	disk[102] = 32'b00110000000000010000000000000001;
	disk[103] = 32'b00110100100000010000000000000100;
	disk[104] = 32'b00101100000000010000000011010110;
	disk[105] = 32'b00001100001001000000000000000000;
	disk[106] = 32'b00110000000000010000000010001000;
	disk[107] = 32'b00110100100000010000000000100111;
	disk[108] = 32'b00101100000000010000000011010110;
	disk[109] = 32'b00001100001001000000000000000000;
	disk[110] = 32'b00110000000000010000000010111101;
	disk[111] = 32'b00110100100000010000000001001010;
	disk[112] = 32'b00101100000000010000000011010110;
	disk[113] = 32'b00001100001001000000000000000000;
	disk[114] = 32'b00110000000000010000000000110100;
	disk[115] = 32'b00110100100000010000000001101101;
	disk[116] = 32'b00101100000000010000000011010110;
	disk[117] = 32'b00001100001001000000000000000000;
	disk[118] = 32'b00110000000000010000000000000001;
	disk[119] = 32'b00110100100000010000000010010000;
	disk[120] = 32'b00101100000000010000000011010110;
	disk[121] = 32'b00001100001001000000000000000000;
	disk[122] = 32'b00110000000000010000000000110110;
	disk[123] = 32'b00110100100000010000000010110011;
	disk[124] = 32'b00101100000000010000000011010110;
	disk[125] = 32'b00001100001001000000000000000000;
	disk[126] = 32'b00110000000000010000000000000001;
	disk[127] = 32'b00001100001000100000000000000000;
	disk[128] = 32'b00001100100000110000000000000000;
	disk[129] = 32'b00001000011000100000100000000000;
	disk[130] = 32'b00110100000000010000000011010110;
	disk[131] = 32'b00101100000000010000000011010110;
	disk[132] = 32'b00001100001001000000000000000000;
	disk[133] = 32'b00110000000000010000000000000001;
	disk[134] = 32'b00110100100000010000000000000100;
	disk[135] = 32'b00101100000000010000000011010110;
	disk[136] = 32'b00001100001001000000000000000000;
	disk[137] = 32'b00110000000000010000000010111110;
	disk[138] = 32'b00110100100000010000000000100111;
	disk[139] = 32'b00101100000000010000000011010110;
	disk[140] = 32'b00001100001001000000000000000000;
	disk[141] = 32'b00110000000000010000000100011001;
	disk[142] = 32'b00110100100000010000000001001010;
	disk[143] = 32'b00101100000000010000000011010110;
	disk[144] = 32'b00001100001001000000000000000000;
	disk[145] = 32'b00110000000000010000000000110101;
	disk[146] = 32'b00110100100000010000000001101101;
	disk[147] = 32'b00101100000000010000000011010110;
	disk[148] = 32'b00001100001001000000000000000000;
	disk[149] = 32'b00110000000000010000000000000001;
	disk[150] = 32'b00110100100000010000000010010000;
	disk[151] = 32'b00101100000000010000000011010110;
	disk[152] = 32'b00001100001001000000000000000000;
	disk[153] = 32'b00110000000000010000000001011100;
	disk[154] = 32'b00110100100000010000000010110011;
	disk[155] = 32'b00101100000000010000000011010110;
	disk[156] = 32'b00001100001001000000000000000000;
	disk[157] = 32'b00110000000000010000000000000001;
	disk[158] = 32'b00001100001000100000000000000000;
	disk[159] = 32'b00001100100000110000000000000000;
	disk[160] = 32'b00001000011000100000100000000000;
	disk[161] = 32'b00110100000000010000000011010110;
	disk[162] = 32'b00101100000000010000000011010110;
	disk[163] = 32'b00001100001001000000000000000000;
	disk[164] = 32'b00110000000000010000000000000001;
	disk[165] = 32'b00110100100000010000000000000100;
	disk[166] = 32'b00101100000000010000000011010110;
	disk[167] = 32'b00001100001001000000000000000000;
	disk[168] = 32'b00110000000000010000000100011010;
	disk[169] = 32'b00110100100000010000000000100111;
	disk[170] = 32'b00101100000000010000000011010110;
	disk[171] = 32'b00001100001001000000000000000000;
	disk[172] = 32'b00110000000000010000000101110111;
	disk[173] = 32'b00110100100000010000000001001010;
	disk[174] = 32'b00101100000000010000000011010110;
	disk[175] = 32'b00001100001001000000000000000000;
	disk[176] = 32'b00110000000000010000000000110110;
	disk[177] = 32'b00110100100000010000000001101101;
	disk[178] = 32'b00101100000000010000000011010110;
	disk[179] = 32'b00001100001001000000000000000000;
	disk[180] = 32'b00110000000000010000000000000001;
	disk[181] = 32'b00110100100000010000000010010000;
	disk[182] = 32'b00101100000000010000000011010110;
	disk[183] = 32'b00001100001001000000000000000000;
	disk[184] = 32'b00110000000000010000000001011110;
	disk[185] = 32'b00110100100000010000000010110011;
	disk[186] = 32'b00101100000000010000000011010110;
	disk[187] = 32'b00001100001001000000000000000000;
	disk[188] = 32'b00110000000000010000000000000001;
	disk[189] = 32'b00001100001000100000000000000000;
	disk[190] = 32'b00001100100000110000000000000000;
	disk[191] = 32'b00001000011000100000100000000000;
	disk[192] = 32'b00110100000000010000000011010110;
	disk[193] = 32'b00101100000000010000000011010110;
	disk[194] = 32'b00001100001001000000000000000000;
	disk[195] = 32'b00110000000000010000000000000001;
	disk[196] = 32'b00110100100000010000000000000100;
	disk[197] = 32'b00101100000000010000000011010110;
	disk[198] = 32'b00001100001001000000000000000000;
	disk[199] = 32'b00110000000000010000000101111000;
	disk[200] = 32'b00110100100000010000000000100111;
	disk[201] = 32'b00101100000000010000000011010110;
	disk[202] = 32'b00001100001001000000000000000000;
	disk[203] = 32'b00110000000000010000000111010101;
	disk[204] = 32'b00110100100000010000000001001010;
	disk[205] = 32'b00101100000000010000000011010110;
	disk[206] = 32'b00001100001001000000000000000000;
	disk[207] = 32'b00110000000000010000000000110111;
	disk[208] = 32'b00110100100000010000000001101101;
	disk[209] = 32'b00101100000000010000000011010110;
	disk[210] = 32'b00001100001001000000000000000000;
	disk[211] = 32'b00110000000000010000000000000001;
	disk[212] = 32'b00110100100000010000000010010000;
	disk[213] = 32'b00101100000000010000000011010110;
	disk[214] = 32'b00001100001001000000000000000000;
	disk[215] = 32'b00110000000000010000000001011110;
	disk[216] = 32'b00110100100000010000000010110011;
	disk[217] = 32'b00101100000000010000000011010110;
	disk[218] = 32'b00001100001001000000000000000000;
	disk[219] = 32'b00110000000000010000000000000001;
	disk[220] = 32'b00001100001000100000000000000000;
	disk[221] = 32'b00001100100000110000000000000000;
	disk[222] = 32'b00001000011000100000100000000000;
	disk[223] = 32'b00110100000000010000000011010110;
	disk[224] = 32'b00101100000000010000000011010110;
	disk[225] = 32'b00001100001001000000000000000000;
	disk[226] = 32'b00110000000000010000000000000001;
	disk[227] = 32'b00110100100000010000000000000100;
	disk[228] = 32'b00101100000000010000000011010110;
	disk[229] = 32'b00001100001001000000000000000000;
	disk[230] = 32'b00110000000000010000000111010110;
	disk[231] = 32'b00110100100000010000000000100111;
	disk[232] = 32'b00101100000000010000000011010110;
	disk[233] = 32'b00001100001001000000000000000000;
	disk[234] = 32'b00110000000000010000001000011110;
	disk[235] = 32'b00110100100000010000000001001010;
	disk[236] = 32'b00101100000000010000000011010110;
	disk[237] = 32'b00001100001001000000000000000000;
	disk[238] = 32'b00110000000000010000000000111000;
	disk[239] = 32'b00110100100000010000000001101101;
	disk[240] = 32'b00101100000000010000000011010110;
	disk[241] = 32'b00001100001001000000000000000000;
	disk[242] = 32'b00110000000000010000000000000001;
	disk[243] = 32'b00110100100000010000000010010000;
	disk[244] = 32'b00101100000000010000000011010110;
	disk[245] = 32'b00001100001001000000000000000000;
	disk[246] = 32'b00110000000000010000000001001001;
	disk[247] = 32'b00110100100000010000000010110011;
	disk[248] = 32'b00101100000000010000000011010110;
	disk[249] = 32'b00001100001001000000000000000000;
	disk[250] = 32'b00110000000000010000000000000001;
	disk[251] = 32'b00001100001000100000000000000000;
	disk[252] = 32'b00001100100000110000000000000000;
	disk[253] = 32'b00001000011000100000100000000000;
	disk[254] = 32'b00110100000000010000000011010110;
	disk[255] = 32'b00101100000000010000000011010110;
	disk[256] = 32'b00001100001001000000000000000000;
	disk[257] = 32'b00110000000000010000000000000001;
	disk[258] = 32'b00110100100000010000000000000100;
	disk[259] = 32'b00101100000000010000000011010110;
	disk[260] = 32'b00001100001001000000000000000000;
	disk[261] = 32'b00110000000000010000001000011111;
	disk[262] = 32'b00110100100000010000000000100111;
	disk[263] = 32'b00101100000000010000000011010110;
	disk[264] = 32'b00001100001001000000000000000000;
	disk[265] = 32'b00110000000000010000001001101001;
	disk[266] = 32'b00110100100000010000000001001010;
	disk[267] = 32'b00101100000000010000000011010110;
	disk[268] = 32'b00001100001001000000000000000000;
	disk[269] = 32'b00110000000000010000000000111001;
	disk[270] = 32'b00110100100000010000000001101101;
	disk[271] = 32'b00101100000000010000000011010110;
	disk[272] = 32'b00001100001001000000000000000000;
	disk[273] = 32'b00110000000000010000000000000001;
	disk[274] = 32'b00110100100000010000000010010000;
	disk[275] = 32'b00101100000000010000000011010110;
	disk[276] = 32'b00001100001001000000000000000000;
	disk[277] = 32'b00110000000000010000000001001011;
	disk[278] = 32'b00110100100000010000000010110011;
	disk[279] = 32'b00101100000000010000000011010110;
	disk[280] = 32'b00001100001001000000000000000000;
	disk[281] = 32'b00110000000000010000000000000001;
	disk[282] = 32'b00001100001000100000000000000000;
	disk[283] = 32'b00001100100000110000000000000000;
	disk[284] = 32'b00001000011000100000100000000000;
	disk[285] = 32'b00110100000000010000000011010110;
	disk[286] = 32'b00101100000000010000000011010110;
	disk[287] = 32'b00001100001001000000000000000000;
	disk[288] = 32'b00110000000000010000000000000001;
	disk[289] = 32'b00110100100000010000000000000100;
	disk[290] = 32'b00101100000000010000000011010110;
	disk[291] = 32'b00001100001001000000000000000000;
	disk[292] = 32'b00110000000000010000001001101010;
	disk[293] = 32'b00110100100000010000000000100111;
	disk[294] = 32'b00101100000000010000000011010110;
	disk[295] = 32'b00001100001001000000000000000000;
	disk[296] = 32'b00110000000000010000001011001000;
	disk[297] = 32'b00110100100000010000000001001010;
	disk[298] = 32'b00101100000000010000000011010110;
	disk[299] = 32'b00001100001001000000000000000000;
	disk[300] = 32'b00110000000000010000000000111010;
	disk[301] = 32'b00110100100000010000000001101101;
	disk[302] = 32'b00101100000000010000000011010110;
	disk[303] = 32'b00001100001001000000000000000000;
	disk[304] = 32'b00110000000000010000000000000001;
	disk[305] = 32'b00110100100000010000000010010000;
	disk[306] = 32'b00101100000000010000000011010110;
	disk[307] = 32'b00001100001001000000000000000000;
	disk[308] = 32'b00110000000000010000000001011111;
	disk[309] = 32'b00110100100000010000000010110011;
	disk[310] = 32'b00101100000000010000000011010110;
	disk[311] = 32'b00001100001001000000000000000000;
	disk[312] = 32'b00110000000000010000000000000001;
	disk[313] = 32'b00001100001000100000000000000000;
	disk[314] = 32'b00001100100000110000000000000000;
	disk[315] = 32'b00001000011000100000100000000000;
	disk[316] = 32'b00110100000000010000000011010110;
	disk[317] = 32'b00101100000000010000000011010110;
	disk[318] = 32'b00001100001001000000000000000000;
	disk[319] = 32'b00110000000000010000000000000001;
	disk[320] = 32'b00110100100000010000000000000100;
	disk[321] = 32'b00101100000000010000000011010110;
	disk[322] = 32'b00001100001001000000000000000000;
	disk[323] = 32'b00110000000000010000001011001001;
	disk[324] = 32'b00110100100000010000000000100111;
	disk[325] = 32'b00101100000000010000000011010110;
	disk[326] = 32'b00001100001001000000000000000000;
	disk[327] = 32'b00110000000000010000001011111000;
	disk[328] = 32'b00110100100000010000000001001010;
	disk[329] = 32'b00101100000000010000000011010110;
	disk[330] = 32'b00001100001001000000000000000000;
	disk[331] = 32'b00110000000000010000000000111011;
	disk[332] = 32'b00110100100000010000000001101101;
	disk[333] = 32'b00101100000000010000000011010110;
	disk[334] = 32'b00001100001001000000000000000000;
	disk[335] = 32'b00110000000000010000000000000001;
	disk[336] = 32'b00110100100000010000000010010000;
	disk[337] = 32'b00101100000000010000000011010110;
	disk[338] = 32'b00001100001001000000000000000000;
	disk[339] = 32'b00110000000000010000000000110000;
	disk[340] = 32'b00110100100000010000000010110011;
	disk[341] = 32'b00101100000000010000000011010110;
	disk[342] = 32'b00001100001001000000000000000000;
	disk[343] = 32'b00110000000000010000000000000001;
	disk[344] = 32'b00001100001000100000000000000000;
	disk[345] = 32'b00001100100000110000000000000000;
	disk[346] = 32'b00001000011000100000100000000000;
	disk[347] = 32'b00110100000000010000000011010110;
	disk[348] = 32'b00111111111000000000000000000000;
	disk[349] = 32'b00110000000000010000000000000001;
	disk[350] = 32'b00110100000000010000000011111011;
	disk[351] = 32'b00110000000000010000000000000010;
	disk[352] = 32'b00110100000000010000000011111100;
	disk[353] = 32'b00110000000000010000000000000011;
	disk[354] = 32'b00110100000000010000000011111101;
	disk[355] = 32'b00110000000000010000000000000100;
	disk[356] = 32'b00110100000000010000000011111110;
	disk[357] = 32'b00110000000000010000000000000101;
	disk[358] = 32'b00110100000000010000000011111111;
	disk[359] = 32'b00110000000000010000000000000110;
	disk[360] = 32'b00110100000000010000000100000000;
	disk[361] = 32'b00110000000000010000000000000111;
	disk[362] = 32'b00110100000000010000000100000001;
	disk[363] = 32'b00110000000000010000000000001000;
	disk[364] = 32'b00110100000000010000000100000010;
	disk[365] = 32'b00110000000000010000000000001001;
	disk[366] = 32'b00110100000000010000000100000011;
	disk[367] = 32'b00110000000000010000000000001010;
	disk[368] = 32'b00110100000000010000000100000100;
	disk[369] = 32'b00110000000000010000000000001011;
	disk[370] = 32'b00110100000000010000000100000101;
	disk[371] = 32'b00110000000000010000000000001100;
	disk[372] = 32'b00110100000000010000000100000110;
	disk[373] = 32'b00110000000000010000000000001101;
	disk[374] = 32'b00110100000000010000000100000111;
	disk[375] = 32'b00110000000000010000000000001110;
	disk[376] = 32'b00110100000000010000000100001000;
	disk[377] = 32'b00110000000000010000000000001111;
	disk[378] = 32'b00110100000000010000000100001001;
	disk[379] = 32'b00110000000000010000011111001111;
	disk[380] = 32'b00110100000000010000000100001010;
	disk[381] = 32'b00110000000000010000000000000101;
	disk[382] = 32'b00110100000000010000000100001011;
	disk[383] = 32'b00101100000000010000000011111011;
	disk[384] = 32'b10011000001000000000000000000000;
	disk[385] = 32'b00001111110111101111111111111111;
	disk[386] = 32'b00110111110111110000000000000000;
	disk[387] = 32'b10000100000000000000000000000010;
	disk[388] = 32'b00101111110111110000000000000000;
	disk[389] = 32'b00001111110111100000000000000001;
	disk[390] = 32'b00111111111000000000000000000000;
	disk[391] = 32'b00111111111000000000000000000000;
	disk[392] = 32'b00110000000000010000000000000000;
	disk[393] = 32'b00110100000000010000000100010001;
	disk[394] = 32'b00101100000000010000000100010001;
	disk[395] = 32'b00001100001001000000000000000000;
	disk[396] = 32'b00101100000000010000000011010110;
	disk[397] = 32'b00001100001000100000000000000000;
	disk[398] = 32'b00001100100000110000000000000000;
	disk[399] = 32'b01110000011000100000000110100010;
	disk[400] = 32'b00101100000000010000000100010001;
	disk[401] = 32'b00101100001000010000000001101101;
	disk[402] = 32'b00001100001001000000000000000000;
	disk[403] = 32'b00101100000000010000000100010000;
	disk[404] = 32'b00001100001000100000000000000000;
	disk[405] = 32'b00001100100000110000000000000000;
	disk[406] = 32'b01011100011000100000000110011010;
	disk[407] = 32'b00101100000000010000000100010001;
	disk[408] = 32'b00001100001111010000000000000000;
	disk[409] = 32'b00111111111000000000000000000000;
	disk[410] = 32'b00101100000000010000000100010001;
	disk[411] = 32'b00001100001001000000000000000000;
	disk[412] = 32'b00110000000000010000000000000001;
	disk[413] = 32'b00001100001000100000000000000000;
	disk[414] = 32'b00001100100000110000000000000000;
	disk[415] = 32'b00001000011000100000100000000000;
	disk[416] = 32'b00110100000000010000000100010001;
	disk[417] = 32'b00111000000000000000000110001010;
	disk[418] = 32'b00110000000000010000000000000000;
	disk[419] = 32'b00001100001111010000000000000000;
	disk[420] = 32'b00111111111000000000000000000000;
	disk[421] = 32'b00110000000000010000000000000000;
	disk[422] = 32'b00110100000000010000000100010011;
	disk[423] = 32'b00110000000000010000000001100011;
	disk[424] = 32'b00110100000000010000000100010100;
	disk[425] = 32'b00101100000000010000000011111111;
	disk[426] = 32'b10011000001000000000000000000000;
	disk[427] = 32'b01111100000000010000000000000000;
	disk[428] = 32'b00110100000000010000000100010101;
	disk[429] = 32'b01111100000000010000000000000000;
	disk[430] = 32'b00110100000000010000000100010110;
	disk[431] = 32'b00101100000000010000000100010011;
	disk[432] = 32'b00001100001001000000000000000000;
	disk[433] = 32'b00101100000000010000000011010110;
	disk[434] = 32'b00001100001000100000000000000000;
	disk[435] = 32'b00001100100000110000000000000000;
	disk[436] = 32'b01110000011000100000000111010010;
	disk[437] = 32'b00101100000000010000000100010011;
	disk[438] = 32'b00101100001000010000000010010000;
	disk[439] = 32'b00001100001001000000000000000000;
	disk[440] = 32'b00110000000000010000000000000000;
	disk[441] = 32'b00001100001000100000000000000000;
	disk[442] = 32'b00001100100000110000000000000000;
	disk[443] = 32'b01011100011000100000000110111111;
	disk[444] = 32'b00110000000000010000000001100011;
	disk[445] = 32'b00110100000000010000000100010011;
	disk[446] = 32'b00111000000000000000000111001010;
	disk[447] = 32'b00101100000000010000000100010011;
	disk[448] = 32'b00101100001000010000000001101101;
	disk[449] = 32'b00001100001001000000000000000000;
	disk[450] = 32'b00101100000000010000000100010101;
	disk[451] = 32'b00001100001000100000000000000000;
	disk[452] = 32'b00001100100000110000000000000000;
	disk[453] = 32'b01011100011000100000000111001010;
	disk[454] = 32'b00101100000000010000000100010011;
	disk[455] = 32'b00110100000000010000000100010100;
	disk[456] = 32'b00110000000000010000000001100011;
	disk[457] = 32'b00110100000000010000000100010011;
	disk[458] = 32'b00101100000000010000000100010011;
	disk[459] = 32'b00001100001001000000000000000000;
	disk[460] = 32'b00110000000000010000000000000001;
	disk[461] = 32'b00001100001000100000000000000000;
	disk[462] = 32'b00001100100000110000000000000000;
	disk[463] = 32'b00001000011000100000100000000000;
	disk[464] = 32'b00110100000000010000000100010011;
	disk[465] = 32'b00111000000000000000000110101111;
	disk[466] = 32'b00101100000000010000000100010100;
	disk[467] = 32'b00001100001001000000000000000000;
	disk[468] = 32'b00101100000000010000000011010110;
	disk[469] = 32'b00001100001000100000000000000000;
	disk[470] = 32'b00001100100000110000000000000000;
	disk[471] = 32'b01110000011000100000000111011101;
	disk[472] = 32'b00101100000000010000000100010100;
	disk[473] = 32'b00001100001001000000000000000000;
	disk[474] = 32'b00101100000000010000000100010110;
	disk[475] = 32'b00110100100000010000000001101101;
	disk[476] = 32'b00111000000000000000000111011111;
	disk[477] = 32'b10000000000000000000000100000111;
	disk[478] = 32'b10000000000000000000000100010101;
	disk[479] = 32'b00111111111000000000000000000000;
	disk[480] = 32'b00101100000000010000000100000000;
	disk[481] = 32'b10011000001000000000000000000000;
	disk[482] = 32'b01111100000000010000000000000000;
	disk[483] = 32'b00110100000000010000000000000011;
	disk[484] = 32'b00101100000000010000000011011000;
	disk[485] = 32'b00110100000000010000000100010111;
	disk[486] = 32'b00110000000000010000000000000001;
	disk[487] = 32'b00110100000000010000000100011000;
	disk[488] = 32'b00101100000000010000000100011000;
	disk[489] = 32'b00001100001001000000000000000000;
	disk[490] = 32'b00110000000000010000000000000000;
	disk[491] = 32'b00001100001000100000000000000000;
	disk[492] = 32'b00001100100000110000000000000000;
	disk[493] = 32'b01100000011000100000001001101101;
	disk[494] = 32'b00101100000000010000000100010111;
	disk[495] = 32'b00101100001000010000000010010000;
	disk[496] = 32'b00001100001001000000000000000000;
	disk[497] = 32'b00110000000000010000000000000000;
	disk[498] = 32'b00001100001000100000000000000000;
	disk[499] = 32'b00001100100000110000000000000000;
	disk[500] = 32'b01011100011000100000000111111011;
	disk[501] = 32'b00110000000000010000000000000000;
	disk[502] = 32'b00110100000000010000000100011000;
	disk[503] = 32'b00101100000000010000000100000111;
	disk[504] = 32'b10011000001000000000000000000000;
	disk[505] = 32'b10000000000000000000000000000011;
	disk[506] = 32'b00111000000000000000001001101100;
	disk[507] = 32'b00101100000000010000000100010111;
	disk[508] = 32'b00101100001000010000000001101101;
	disk[509] = 32'b00001100001001000000000000000000;
	disk[510] = 32'b00101100000000010000000000000011;
	disk[511] = 32'b00001100001000100000000000000000;
	disk[512] = 32'b00001100100000110000000000000000;
	disk[513] = 32'b01011100011000100000001001100101;
	disk[514] = 32'b00101100000000010000000100010111;
	disk[515] = 32'b00001100001001000000000000000000;
	disk[516] = 32'b00110000000000010000000000000000;
	disk[517] = 32'b00110100100000010000000010010000;
	disk[518] = 32'b00110000000000010000000000000000;
	disk[519] = 32'b00110100000000010000000100011000;
	disk[520] = 32'b00101100000000010000000011010110;
	disk[521] = 32'b00001100001001000000000000000000;
	disk[522] = 32'b00101100000000010000000100010111;
	disk[523] = 32'b00001100001000100000000000000000;
	disk[524] = 32'b00001100100000110000000000000000;
	disk[525] = 32'b01100000011000100000001001100101;
	disk[526] = 32'b00101100000000010000000100010111;
	disk[527] = 32'b00001100001001000000000000000000;
	disk[528] = 32'b00110000000000010000000000000001;
	disk[529] = 32'b00001100001000100000000000000000;
	disk[530] = 32'b00001100100000110000000000000000;
	disk[531] = 32'b00001000011000100000100000000000;
	disk[532] = 32'b00101100001000010000000010010000;
	disk[533] = 32'b00001100001001000000000000000000;
	disk[534] = 32'b00110000000000010000000000000000;
	disk[535] = 32'b00001100001000100000000000000000;
	disk[536] = 32'b00001100100000110000000000000000;
	disk[537] = 32'b01100000011000100000001001011110;
	disk[538] = 32'b00101100000000010000000100010111;
	disk[539] = 32'b00001100001001000000000000000000;
	disk[540] = 32'b00101100000000010000000100010111;
	disk[541] = 32'b00001100001001010000000000000000;
	disk[542] = 32'b00110000000000010000000000000001;
	disk[543] = 32'b00001100001000100000000000000000;
	disk[544] = 32'b00001100101000110000000000000000;
	disk[545] = 32'b00001000011000100000100000000000;
	disk[546] = 32'b00101100001000010000000000000100;
	disk[547] = 32'b00110100100000010000000000000100;
	disk[548] = 32'b00101100000000010000000100010111;
	disk[549] = 32'b00001100001001000000000000000000;
	disk[550] = 32'b00101100000000010000000100010111;
	disk[551] = 32'b00001100001001010000000000000000;
	disk[552] = 32'b00110000000000010000000000000001;
	disk[553] = 32'b00001100001000100000000000000000;
	disk[554] = 32'b00001100101000110000000000000000;
	disk[555] = 32'b00001000011000100000100000000000;
	disk[556] = 32'b00101100001000010000000000100111;
	disk[557] = 32'b00110100100000010000000000100111;
	disk[558] = 32'b00101100000000010000000100010111;
	disk[559] = 32'b00001100001001000000000000000000;
	disk[560] = 32'b00101100000000010000000100010111;
	disk[561] = 32'b00001100001001010000000000000000;
	disk[562] = 32'b00110000000000010000000000000001;
	disk[563] = 32'b00001100001000100000000000000000;
	disk[564] = 32'b00001100101000110000000000000000;
	disk[565] = 32'b00001000011000100000100000000000;
	disk[566] = 32'b00101100001000010000000001001010;
	disk[567] = 32'b00110100100000010000000001001010;
	disk[568] = 32'b00101100000000010000000100010111;
	disk[569] = 32'b00001100001001000000000000000000;
	disk[570] = 32'b00101100000000010000000100010111;
	disk[571] = 32'b00001100001001010000000000000000;
	disk[572] = 32'b00110000000000010000000000000001;
	disk[573] = 32'b00001100001000100000000000000000;
	disk[574] = 32'b00001100101000110000000000000000;
	disk[575] = 32'b00001000011000100000100000000000;
	disk[576] = 32'b00101100001000010000000001101101;
	disk[577] = 32'b00110100100000010000000001101101;
	disk[578] = 32'b00101100000000010000000100010111;
	disk[579] = 32'b00001100001001000000000000000000;
	disk[580] = 32'b00101100000000010000000100010111;
	disk[581] = 32'b00001100001001010000000000000000;
	disk[582] = 32'b00110000000000010000000000000001;
	disk[583] = 32'b00001100001000100000000000000000;
	disk[584] = 32'b00001100101000110000000000000000;
	disk[585] = 32'b00001000011000100000100000000000;
	disk[586] = 32'b00101100001000010000000010010000;
	disk[587] = 32'b00110100100000010000000010010000;
	disk[588] = 32'b00101100000000010000000100010111;
	disk[589] = 32'b00001100001001000000000000000000;
	disk[590] = 32'b00101100000000010000000100010111;
	disk[591] = 32'b00001100001001010000000000000000;
	disk[592] = 32'b00110000000000010000000000000001;
	disk[593] = 32'b00001100001000100000000000000000;
	disk[594] = 32'b00001100101000110000000000000000;
	disk[595] = 32'b00001000011000100000100000000000;
	disk[596] = 32'b00101100001000010000000010110011;
	disk[597] = 32'b00110100100000010000000010110011;
	disk[598] = 32'b00101100000000010000000100010111;
	disk[599] = 32'b00001100001001000000000000000000;
	disk[600] = 32'b00110000000000010000000000000001;
	disk[601] = 32'b00001100001000100000000000000000;
	disk[602] = 32'b00001100100000110000000000000000;
	disk[603] = 32'b00001000011000100000100000000000;
	disk[604] = 32'b00110100000000010000000100010111;
	disk[605] = 32'b00111000000000000000001000001110;
	disk[606] = 32'b00101100000000010000000011010110;
	disk[607] = 32'b00001100001001000000000000000000;
	disk[608] = 32'b00110000000000010000000000000001;
	disk[609] = 32'b00001100001000100000000000000000;
	disk[610] = 32'b00001100100000110000000000000000;
	disk[611] = 32'b00010000011000100000100000000000;
	disk[612] = 32'b00110100000000010000000011010110;
	disk[613] = 32'b00101100000000010000000100010111;
	disk[614] = 32'b00001100001001000000000000000000;
	disk[615] = 32'b00110000000000010000000000000001;
	disk[616] = 32'b00001100001000100000000000000000;
	disk[617] = 32'b00001100100000110000000000000000;
	disk[618] = 32'b00001000011000100000100000000000;
	disk[619] = 32'b00110100000000010000000100010111;
	disk[620] = 32'b00111000000000000000000111101000;
	disk[621] = 32'b00111111111000000000000000000000;
	disk[622] = 32'b00110000000000010000000000000000;
	disk[623] = 32'b00110100000000010000000100011111;
	disk[624] = 32'b00110000000000010000000000000000;
	disk[625] = 32'b00110100000000010000000100011101;
	disk[626] = 32'b00110000000000010000000000000000;
	disk[627] = 32'b00110100000000010000000100011110;
	disk[628] = 32'b00101100000000010000000011010110;
	disk[629] = 32'b00001100001001000000000000000000;
	disk[630] = 32'b00110000000000010000000000000001;
	disk[631] = 32'b00001100001000100000000000000000;
	disk[632] = 32'b00001100100000110000000000000000;
	disk[633] = 32'b00010000011000100000100000000000;
	disk[634] = 32'b00101100001000010000000001001010;
	disk[635] = 32'b00110100000000010000000100100000;
	disk[636] = 32'b00101100000000010000000011010111;
	disk[637] = 32'b00110100000000010000000100100001;
	disk[638] = 32'b00110000000000010000000000000000;
	disk[639] = 32'b00110100000000010000000100011111;
	disk[640] = 32'b00101100000000010000000011111100;
	disk[641] = 32'b10011000001000000000000000000000;
	disk[642] = 32'b01111100000000010000000000000000;
	disk[643] = 32'b00110100000000010000000100011011;
	disk[644] = 32'b00001111110111101111111111111111;
	disk[645] = 32'b00110111110111110000000000000000;
	disk[646] = 32'b00101100000000010000000100011011;
	disk[647] = 32'b00110100000000010000000101011011;
	disk[648] = 32'b00101100000000010000000101011011;
	disk[649] = 32'b00110100000000010000000100010000;
	disk[650] = 32'b10000100000000000000000110001000;
	disk[651] = 32'b00101111110111110000000000000000;
	disk[652] = 32'b00001111110111100000000000000001;
	disk[653] = 32'b00001111101000010000000000000000;
	disk[654] = 32'b00110100000000010000000100011100;
	disk[655] = 32'b00101100000000010000000100011100;
	disk[656] = 32'b00001100001001000000000000000000;
	disk[657] = 32'b00110000000000010000000000000000;
	disk[658] = 32'b00001100001000100000000000000000;
	disk[659] = 32'b00001100100000110000000000000000;
	disk[660] = 32'b01100000011000100000001010011001;
	disk[661] = 32'b00101100000000010000000100001000;
	disk[662] = 32'b10011000001000000000000000000000;
	disk[663] = 32'b10000000000000000000000100011011;
	disk[664] = 32'b00111111111000000000000000000000;
	disk[665] = 32'b00101100000000010000000100011111;
	disk[666] = 32'b00001100001001000000000000000000;
	disk[667] = 32'b00110000000000010000000000000000;
	disk[668] = 32'b00001100001001010000000000000000;
	disk[669] = 32'b00110000000000010000000000000001;
	disk[670] = 32'b00001100001000100000000000000000;
	disk[671] = 32'b00001100101000110000000000000000;
	disk[672] = 32'b00010000011000100000100000000000;
	disk[673] = 32'b00001100001000100000000000000000;
	disk[674] = 32'b00001100100000110000000000000000;
	disk[675] = 32'b01100000011000100000001011011101;
	disk[676] = 32'b00101100000000010000000011111101;
	disk[677] = 32'b10011000001000000000000000000000;
	disk[678] = 32'b01111100000000010000000000000000;
	disk[679] = 32'b00110100000000010000000100011101;
	disk[680] = 32'b01111100000000010000000000000000;
	disk[681] = 32'b00110100000000010000000100011110;
	disk[682] = 32'b00101100000000010000000100011101;
	disk[683] = 32'b00001100001101000000000000000000;
	disk[684] = 32'b00101100000000010000000100011110;
	disk[685] = 32'b00001100001101010000000000000000;
	disk[686] = 32'b00101010101101010000010000000000;
	disk[687] = 32'b01001010100101010000100000000000;
	disk[688] = 32'b00001100001111010000000000000000;
	disk[689] = 32'b00110100000000010000000100011010;
	disk[690] = 32'b00101100000000010000000100100000;
	disk[691] = 32'b00001100001001000000000000000000;
	disk[692] = 32'b00101100000000010000000100001010;
	disk[693] = 32'b00001100001000100000000000000000;
	disk[694] = 32'b00001100100000110000000000000000;
	disk[695] = 32'b01011100011000100000001011000010;
	disk[696] = 32'b00110000000000010000000000000000;
	disk[697] = 32'b00110100000000010000000100100000;
	disk[698] = 32'b00101100000000010000000100100001;
	disk[699] = 32'b00001100001001000000000000000000;
	disk[700] = 32'b00110000000000010000000000000001;
	disk[701] = 32'b00001100001000100000000000000000;
	disk[702] = 32'b00001100100000110000000000000000;
	disk[703] = 32'b00001000011000100000100000000000;
	disk[704] = 32'b00110100000000010000000100100001;
	disk[705] = 32'b00111000000000000000001011001001;
	disk[706] = 32'b00101100000000010000000100100000;
	disk[707] = 32'b00001100001001000000000000000000;
	disk[708] = 32'b00110000000000010000000000000001;
	disk[709] = 32'b00001100001000100000000000000000;
	disk[710] = 32'b00001100100000110000000000000000;
	disk[711] = 32'b00001000011000100000100000000000;
	disk[712] = 32'b00110100000000010000000100100000;
	disk[713] = 32'b00101100000000010000000100011010;
	disk[714] = 32'b10110100000000010000000000000000;
	disk[715] = 32'b00101100000000010000000100100001;
	disk[716] = 32'b00001100001000100000000000000000;
	disk[717] = 32'b00101100000000010000000100100000;
	disk[718] = 32'b00001100001000110000000000000000;
	disk[719] = 32'b10011100011000100000000000000000;
	disk[720] = 32'b00101100000000010000000100011001;
	disk[721] = 32'b00001100001001000000000000000000;
	disk[722] = 32'b00110000000000010000000000000001;
	disk[723] = 32'b00001100001000100000000000000000;
	disk[724] = 32'b00001100100000110000000000000000;
	disk[725] = 32'b00001000011000100000100000000000;
	disk[726] = 32'b00110100000000010000000100011001;
	disk[727] = 32'b10000000000000000000000100011001;
	disk[728] = 32'b00101100000000010000000011111110;
	disk[729] = 32'b10011000001000000000000000000000;
	disk[730] = 32'b01111100000000010000000000000000;
	disk[731] = 32'b00110100000000010000000100011111;
	disk[732] = 32'b00111000000000000000001010011001;
	disk[733] = 32'b00101100000000010000000100011001;
	disk[734] = 32'b00001100001001000000000000000000;
	disk[735] = 32'b00110000000000010000000000000000;
	disk[736] = 32'b00001100001000100000000000000000;
	disk[737] = 32'b00001100100000110000000000000000;
	disk[738] = 32'b01100000011000100000001100011110;
	disk[739] = 32'b00101100000000010000000100000110;
	disk[740] = 32'b10011000001000000000000000000000;
	disk[741] = 32'b01111100000000010000000000000000;
	disk[742] = 32'b00110100000000010000000100011111;
	disk[743] = 32'b00101100000000010000000100011111;
	disk[744] = 32'b00001100001001000000000000000000;
	disk[745] = 32'b00110000000000010000000000000001;
	disk[746] = 32'b00001100001000100000000000000000;
	disk[747] = 32'b00001100100000110000000000000000;
	disk[748] = 32'b01011100011000100000001100011110;
	disk[749] = 32'b00101100000000010000000011010110;
	disk[750] = 32'b00001100001001000000000000000000;
	disk[751] = 32'b00101100000000010000000011010111;
	disk[752] = 32'b00110100100000010000000000000100;
	disk[753] = 32'b00101100000000010000000011010110;
	disk[754] = 32'b00001100001001000000000000000000;
	disk[755] = 32'b00101100000000010000000011010110;
	disk[756] = 32'b00001100001001010000000000000000;
	disk[757] = 32'b00110000000000010000000000000001;
	disk[758] = 32'b00001100001000100000000000000000;
	disk[759] = 32'b00001100101000110000000000000000;
	disk[760] = 32'b00010000011000100000100000000000;
	disk[761] = 32'b00101100001000010000000001001010;
	disk[762] = 32'b00001100001001010000000000000000;
	disk[763] = 32'b00110000000000010000000000000001;
	disk[764] = 32'b00001100001000100000000000000000;
	disk[765] = 32'b00001100101000110000000000000000;
	disk[766] = 32'b00001000011000100000100000000000;
	disk[767] = 32'b00110100100000010000000000100111;
	disk[768] = 32'b00101100000000010000000011010110;
	disk[769] = 32'b00001100001001000000000000000000;
	disk[770] = 32'b00101100000000010000000100100000;
	disk[771] = 32'b00001100001001010000000000000000;
	disk[772] = 32'b00110000000000010000000000000001;
	disk[773] = 32'b00001100001000100000000000000000;
	disk[774] = 32'b00001100101000110000000000000000;
	disk[775] = 32'b00010000011000100000100000000000;
	disk[776] = 32'b00110100100000010000000001001010;
	disk[777] = 32'b00101100000000010000000011010110;
	disk[778] = 32'b00001100001001000000000000000000;
	disk[779] = 32'b00101100000000010000000100011011;
	disk[780] = 32'b00110100100000010000000001101101;
	disk[781] = 32'b00101100000000010000000011010110;
	disk[782] = 32'b00001100001001000000000000000000;
	disk[783] = 32'b00110000000000010000000000000001;
	disk[784] = 32'b00110100100000010000000010010000;
	disk[785] = 32'b00101100000000010000000011010110;
	disk[786] = 32'b00001100001001000000000000000000;
	disk[787] = 32'b00101100000000010000000100011001;
	disk[788] = 32'b00110100100000010000000010110011;
	disk[789] = 32'b00101100000000010000000011010110;
	disk[790] = 32'b00001100001001000000000000000000;
	disk[791] = 32'b00110000000000010000000000000001;
	disk[792] = 32'b00001100001000100000000000000000;
	disk[793] = 32'b00001100100000110000000000000000;
	disk[794] = 32'b00001000011000100000100000000000;
	disk[795] = 32'b00110100000000010000000011010110;
	disk[796] = 32'b00101100000000010000000100100001;
	disk[797] = 32'b00110100000000010000000011010111;
	disk[798] = 32'b00111111111000000000000000000000;
	disk[799] = 32'b01111100000000010000000000000000;
	disk[800] = 32'b00110100000000010000000100100010;
	disk[801] = 32'b00101100000000010000000100100010;
	disk[802] = 32'b10110100000000010000000000000000;
	disk[803] = 32'b00111111111000000000000000000000;
	disk[804] = 32'b10110000000000010000000000000000;
	disk[805] = 32'b00110100000000010000000100100011;
	disk[806] = 32'b10000000000000000000000100100011;
	disk[807] = 32'b00111111111000000000000000000000;
	disk[808] = 32'b00001111110111101111111111111111;
	disk[809] = 32'b00110111110111110000000000000000;
	disk[810] = 32'b00101100000000010000000100100100;
	disk[811] = 32'b00110100000000010000000101011011;
	disk[812] = 32'b00101100000000010000000101011011;
	disk[813] = 32'b00110100000000010000000100010000;
	disk[814] = 32'b10000100000000000000000110001000;
	disk[815] = 32'b00101111110111110000000000000000;
	disk[816] = 32'b00001111110111100000000000000001;
	disk[817] = 32'b00001111101000010000000000000000;
	disk[818] = 32'b00110100000000010000000100100101;
	disk[819] = 32'b00101100000000010000000100100101;
	disk[820] = 32'b00001100001001000000000000000000;
	disk[821] = 32'b00110000000000010000000000000000;
	disk[822] = 32'b00001100001000100000000000000000;
	disk[823] = 32'b00001100100000110000000000000000;
	disk[824] = 32'b01100000011000100000001101110000;
	disk[825] = 32'b00110000000000010000000000000000;
	disk[826] = 32'b00110100000000010000000100101000;
	disk[827] = 32'b00101100000000010000000100100101;
	disk[828] = 32'b00101100001000010000000000100111;
	disk[829] = 32'b00110100000000010000000100100110;
	disk[830] = 32'b00101100000000010000000100100101;
	disk[831] = 32'b00101100001000010000000000000100;
	disk[832] = 32'b00110100000000010000000100100111;
	disk[833] = 32'b00000000000000000000000000000000;
	disk[834] = 32'b00101100000000010000000100101000;
	disk[835] = 32'b00001100001001000000000000000000;
	disk[836] = 32'b00101100000000010000000100100101;
	disk[837] = 32'b00101100001000010000000010110011;
	disk[838] = 32'b00001100001000100000000000000000;
	disk[839] = 32'b00001100100000110000000000000000;
	disk[840] = 32'b01110000011000100000001101110000;
	disk[841] = 32'b00101100000000010000000100100111;
	disk[842] = 32'b00001100001000100000000000000000;
	disk[843] = 32'b00101100000000010000000100100110;
	disk[844] = 32'b00001100001000110000000000000000;
	disk[845] = 32'b00110000000000010000000000000001;
	disk[846] = 32'b10010100000000010000000000000000;
	disk[847] = 32'b10001000011000100000000000000000;
	disk[848] = 32'b10010100000000000000000000000000;
	disk[849] = 32'b00101100000000010000000100100110;
	disk[850] = 32'b00001100001001000000000000000000;
	disk[851] = 32'b00101100000000010000000100001010;
	disk[852] = 32'b00001100001000100000000000000000;
	disk[853] = 32'b00001100100000110000000000000000;
	disk[854] = 32'b01011100011000100000001101100001;
	disk[855] = 32'b00110000000000010000000000000000;
	disk[856] = 32'b00110100000000010000000100100110;
	disk[857] = 32'b00101100000000010000000100100111;
	disk[858] = 32'b00001100001001000000000000000000;
	disk[859] = 32'b00110000000000010000000000000001;
	disk[860] = 32'b00001100001000100000000000000000;
	disk[861] = 32'b00001100100000110000000000000000;
	disk[862] = 32'b00001000011000100000100000000000;
	disk[863] = 32'b00110100000000010000000100100111;
	disk[864] = 32'b00111000000000000000001101101000;
	disk[865] = 32'b00101100000000010000000100100110;
	disk[866] = 32'b00001100001001000000000000000000;
	disk[867] = 32'b00110000000000010000000000000001;
	disk[868] = 32'b00001100001000100000000000000000;
	disk[869] = 32'b00001100100000110000000000000000;
	disk[870] = 32'b00001000011000100000100000000000;
	disk[871] = 32'b00110100000000010000000100100110;
	disk[872] = 32'b00101100000000010000000100101000;
	disk[873] = 32'b00001100001001000000000000000000;
	disk[874] = 32'b00110000000000010000000000000001;
	disk[875] = 32'b00001100001000100000000000000000;
	disk[876] = 32'b00001100100000110000000000000000;
	disk[877] = 32'b00001000011000100000100000000000;
	disk[878] = 32'b00110100000000010000000100101000;
	disk[879] = 32'b00111000000000000000001101000010;
	disk[880] = 32'b00111111111000000000000000000000;
	disk[881] = 32'b00101100000000010000000100101001;
	disk[882] = 32'b00001100001110100000000000000000;
	disk[883] = 32'b00110000000110110000000000100000;
	disk[884] = 32'b00011011010110111101100000000000;
	disk[885] = 32'b00001111010110100000000000000001;
	disk[886] = 32'b11000111011000010000000101011110;
	disk[887] = 32'b00001111011110110000000000000001;
	disk[888] = 32'b11000111011000100000000101011110;
	disk[889] = 32'b00001111011110110000000000000001;
	disk[890] = 32'b11000111011000110000000101011110;
	disk[891] = 32'b00001111011110110000000000000001;
	disk[892] = 32'b11000111011001000000000101011110;
	disk[893] = 32'b00001111011110110000000000000001;
	disk[894] = 32'b11000111011001010000000101011110;
	disk[895] = 32'b00001111011110110000000000000001;
	disk[896] = 32'b11000111011111010000000101011110;
	disk[897] = 32'b00001111011110110000000000000001;
	disk[898] = 32'b11000111011111100000000101011110;
	disk[899] = 32'b00001111011110110000000000000001;
	disk[900] = 32'b11000111011111110000000101011110;
	disk[901] = 32'b00001111011110110000000000000001;
	disk[902] = 32'b00111111111000000000000000000000;
	disk[903] = 32'b00101100000000010000000100101010;
	disk[904] = 32'b00001100001110100000000000000000;
	disk[905] = 32'b00110000000110110000000000100000;
	disk[906] = 32'b00011011010110111101100000000000;
	disk[907] = 32'b00001111010110100000000000000001;
	disk[908] = 32'b11001011011000010000000101011110;
	disk[909] = 32'b00001111011110110000000000000001;
	disk[910] = 32'b11001011011000100000000101011110;
	disk[911] = 32'b00001111011110110000000000000001;
	disk[912] = 32'b11001011011000110000000101011110;
	disk[913] = 32'b00001111011110110000000000000001;
	disk[914] = 32'b11001011011001000000000101011110;
	disk[915] = 32'b00001111011110110000000000000001;
	disk[916] = 32'b11001011011001010000000101011110;
	disk[917] = 32'b00001111011110110000000000000001;
	disk[918] = 32'b11001011011111010000000101011110;
	disk[919] = 32'b00001111011110110000000000000001;
	disk[920] = 32'b11001011011111100000000101011110;
	disk[921] = 32'b00001111011110110000000000000001;
	disk[922] = 32'b11001011011111110000000101011110;
	disk[923] = 32'b00001111011110110000000000000001;
	disk[924] = 32'b00111111111000000000000000000000;
	disk[925] = 32'b00110000000000010000000000000000;
	disk[926] = 32'b00110100000000010000000100101100;
	disk[927] = 32'b00101100000000010000000100000001;
	disk[928] = 32'b10011000001000000000000000000000;
	disk[929] = 32'b01111100000000010000000000000000;
	disk[930] = 32'b00110100000000010000000100001100;
	disk[931] = 32'b00101100000000010000000100101100;
	disk[932] = 32'b00001100001001000000000000000000;
	disk[933] = 32'b00101100000000010000000100001100;
	disk[934] = 32'b00001100001000100000000000000000;
	disk[935] = 32'b00001100100000110000000000000000;
	disk[936] = 32'b01110000011000100000001111011100;
	disk[937] = 32'b00101100000000010000000100000011;
	disk[938] = 32'b10011000001000000000000000000000;
	disk[939] = 32'b10000000000000000000000100101100;
	disk[940] = 32'b01111100000000010000000000000000;
	disk[941] = 32'b00110100000000010000000100101011;
	disk[942] = 32'b00001111110111101111111111111111;
	disk[943] = 32'b00110111110111110000000000000000;
	disk[944] = 32'b00101100000000010000000100101011;
	disk[945] = 32'b00110100000000010000000101011011;
	disk[946] = 32'b00101100000000010000000101011011;
	disk[947] = 32'b00110100000000010000000100010000;
	disk[948] = 32'b10000100000000000000000110001000;
	disk[949] = 32'b00101111110111110000000000000000;
	disk[950] = 32'b00001111110111100000000000000001;
	disk[951] = 32'b00001111101000010000000000000000;
	disk[952] = 32'b00110100000000010000000100101101;
	disk[953] = 32'b00101100000000010000000100101101;
	disk[954] = 32'b00001100001001000000000000000000;
	disk[955] = 32'b00110000000000010000000000000000;
	disk[956] = 32'b00001100001000100000000000000000;
	disk[957] = 32'b00001100100000110000000000000000;
	disk[958] = 32'b01100000011000100000001111011000;
	disk[959] = 32'b00101100000000010000000100101100;
	disk[960] = 32'b00001100001001000000000000000000;
	disk[961] = 32'b00101100000000010000000100101011;
	disk[962] = 32'b00110100100000010000000011011001;
	disk[963] = 32'b00101100000000010000000100101100;
	disk[964] = 32'b00001100001001000000000000000000;
	disk[965] = 32'b00101100000000010000000100101100;
	disk[966] = 32'b00001100001001010000000000000000;
	disk[967] = 32'b00110000000000010000000000000001;
	disk[968] = 32'b00001100001000100000000000000000;
	disk[969] = 32'b00001100101000110000000000000000;
	disk[970] = 32'b00001000011000100000100000000000;
	disk[971] = 32'b00110100100000010000000011100011;
	disk[972] = 32'b00101100000000010000000100101100;
	disk[973] = 32'b00001100001001000000000000000000;
	disk[974] = 32'b00110000000000010000000000000000;
	disk[975] = 32'b00110100100000010000000011101101;
	disk[976] = 32'b00101100000000010000000100101100;
	disk[977] = 32'b00001100001001000000000000000000;
	disk[978] = 32'b00110000000000010000000000000001;
	disk[979] = 32'b00001100001000100000000000000000;
	disk[980] = 32'b00001100100000110000000000000000;
	disk[981] = 32'b00001000011000100000100000000000;
	disk[982] = 32'b00110100000000010000000100101100;
	disk[983] = 32'b00111000000000000000001111011011;
	disk[984] = 32'b00101100000000010000000100000111;
	disk[985] = 32'b10011000001000000000000000000000;
	disk[986] = 32'b10000000000000000000000100101011;
	disk[987] = 32'b00111000000000000000001110100011;
	disk[988] = 32'b00101100000000010000000100101100;
	disk[989] = 32'b00001100001001000000000000000000;
	disk[990] = 32'b00110000000000010000000000001010;
	disk[991] = 32'b00001100001000100000000000000000;
	disk[992] = 32'b00001100100000110000000000000000;
	disk[993] = 32'b01110000011000100000001111110110;
	disk[994] = 32'b00101100000000010000000100101100;
	disk[995] = 32'b00001100001001000000000000000000;
	disk[996] = 32'b00110000000000010000000000000000;
	disk[997] = 32'b00110100100000010000000011011001;
	disk[998] = 32'b00101100000000010000000100101100;
	disk[999] = 32'b00001100001001000000000000000000;
	disk[1000] = 32'b00110000000000010000000000000000;
	disk[1001] = 32'b00110100100000010000000011100011;
	disk[1002] = 32'b00101100000000010000000100101100;
	disk[1003] = 32'b00001100001001000000000000000000;
	disk[1004] = 32'b00110000000000010000000000000000;
	disk[1005] = 32'b00110100100000010000000011101101;
	disk[1006] = 32'b00101100000000010000000100101100;
	disk[1007] = 32'b00001100001001000000000000000000;
	disk[1008] = 32'b00110000000000010000000000000001;
	disk[1009] = 32'b00001100001000100000000000000000;
	disk[1010] = 32'b00001100100000110000000000000000;
	disk[1011] = 32'b00001000011000100000100000000000;
	disk[1012] = 32'b00110100000000010000000100101100;
	disk[1013] = 32'b00111000000000000000001111011100;
	disk[1014] = 32'b00101100000000010000000100000010;
	disk[1015] = 32'b10011000001000000000000000000000;
	disk[1016] = 32'b00111111111000000000000000000000;
	disk[1017] = 32'b00110000000000010000000000000000;
	disk[1018] = 32'b00110100000000010000000100101110;
	disk[1019] = 32'b00110000000000010000000000000001;
	disk[1020] = 32'b00110100000000010000000100110001;
	disk[1021] = 32'b00110000000000010000000000000000;
	disk[1022] = 32'b00110100000000010000000100110011;
	disk[1023] = 32'b00001111110111101111111111111111;
	disk[1024] = 32'b00110111110111110000000000000000;
	disk[1025] = 32'b10000100000000000000001110011101;
	disk[1026] = 32'b00101111110111110000000000000000;
	disk[1027] = 32'b00001111110111100000000000000001;
	disk[1028] = 32'b00101100000000010000000100001001;
	disk[1029] = 32'b10011000001000000000000000000000;
	disk[1030] = 32'b01111100000000010000000000000000;
	disk[1031] = 32'b00110100000000010000000100101111;
	disk[1032] = 32'b00101100000000010000000100101111;
	disk[1033] = 32'b10111100000000010000000000000000;
	disk[1034] = 32'b00101100000000010000000100001100;
	disk[1035] = 32'b00110100000000010000000100110000;
	disk[1036] = 32'b00110000000000010000000000000000;
	disk[1037] = 32'b10100100001000000000000000000000;
	disk[1038] = 32'b00101100000000010000000100110000;
	disk[1039] = 32'b00001100001001000000000000000000;
	disk[1040] = 32'b00110000000000010000000000000000;
	disk[1041] = 32'b00001100001000100000000000000000;
	disk[1042] = 32'b00001100100000110000000000000000;
	disk[1043] = 32'b01101100011000100000010100110001;
	disk[1044] = 32'b00101100000000010000000100110001;
	disk[1045] = 32'b00001100001001000000000000000000;
	disk[1046] = 32'b00110000000000010000000000000000;
	disk[1047] = 32'b00001100001000100000000000000000;
	disk[1048] = 32'b00001100100000110000000000000000;
	disk[1049] = 32'b01100000011000100000010010111001;
	disk[1050] = 32'b00101100000000010000000100110011;
	disk[1051] = 32'b00001100001001000000000000000000;
	disk[1052] = 32'b00110000000000010000000000000001;
	disk[1053] = 32'b00001100001000100000000000000000;
	disk[1054] = 32'b00001100100000110000000000000000;
	disk[1055] = 32'b01011100011000100000010001110011;
	disk[1056] = 32'b00101100000000010000000100101110;
	disk[1057] = 32'b00001100001001000000000000000000;
	disk[1058] = 32'b00101100000000010000000100110000;
	disk[1059] = 32'b00001100001001010000000000000000;
	disk[1060] = 32'b00110000000000010000000000000001;
	disk[1061] = 32'b00001100001000100000000000000000;
	disk[1062] = 32'b00001100101000110000000000000000;
	disk[1063] = 32'b00010000011000100000100000000000;
	disk[1064] = 32'b00001100001000100000000000000000;
	disk[1065] = 32'b00001100100000110000000000000000;
	disk[1066] = 32'b01110000011000100000010001011110;
	disk[1067] = 32'b00101100000000010000000100101110;
	disk[1068] = 32'b00110100000000010000000100110010;
	disk[1069] = 32'b00101100000000010000000100110010;
	disk[1070] = 32'b00001100001001000000000000000000;
	disk[1071] = 32'b00101100000000010000000100110000;
	disk[1072] = 32'b00001100001001010000000000000000;
	disk[1073] = 32'b00110000000000010000000000000001;
	disk[1074] = 32'b00001100001000100000000000000000;
	disk[1075] = 32'b00001100101000110000000000000000;
	disk[1076] = 32'b00010000011000100000100000000000;
	disk[1077] = 32'b00001100001000100000000000000000;
	disk[1078] = 32'b00001100100000110000000000000000;
	disk[1079] = 32'b01110000011000100000010001011110;
	disk[1080] = 32'b00101100000000010000000100110010;
	disk[1081] = 32'b00001100001001000000000000000000;
	disk[1082] = 32'b00101100000000010000000100110010;
	disk[1083] = 32'b00001100001001010000000000000000;
	disk[1084] = 32'b00110000000000010000000000000001;
	disk[1085] = 32'b00001100001000100000000000000000;
	disk[1086] = 32'b00001100101000110000000000000000;
	disk[1087] = 32'b00001000011000100000100000000000;
	disk[1088] = 32'b00101100001000010000000011101101;
	disk[1089] = 32'b00110100100000010000000011101101;
	disk[1090] = 32'b00101100000000010000000100110010;
	disk[1091] = 32'b00001100001001000000000000000000;
	disk[1092] = 32'b00101100000000010000000100110010;
	disk[1093] = 32'b00001100001001010000000000000000;
	disk[1094] = 32'b00110000000000010000000000000001;
	disk[1095] = 32'b00001100001000100000000000000000;
	disk[1096] = 32'b00001100101000110000000000000000;
	disk[1097] = 32'b00001000011000100000100000000000;
	disk[1098] = 32'b00101100001000010000000011011001;
	disk[1099] = 32'b00110100100000010000000011011001;
	disk[1100] = 32'b00101100000000010000000100110010;
	disk[1101] = 32'b00001100001001000000000000000000;
	disk[1102] = 32'b00101100000000010000000100110010;
	disk[1103] = 32'b00001100001001010000000000000000;
	disk[1104] = 32'b00110000000000010000000000000001;
	disk[1105] = 32'b00001100001000100000000000000000;
	disk[1106] = 32'b00001100101000110000000000000000;
	disk[1107] = 32'b00001000011000100000100000000000;
	disk[1108] = 32'b00101100001000010000000011100011;
	disk[1109] = 32'b00110100100000010000000011100011;
	disk[1110] = 32'b00101100000000010000000100110010;
	disk[1111] = 32'b00001100001001000000000000000000;
	disk[1112] = 32'b00110000000000010000000000000001;
	disk[1113] = 32'b00001100001000100000000000000000;
	disk[1114] = 32'b00001100100000110000000000000000;
	disk[1115] = 32'b00001000011000100000100000000000;
	disk[1116] = 32'b00110100000000010000000100110010;
	disk[1117] = 32'b00111000000000000000010000101101;
	disk[1118] = 32'b00101100000000010000000100101110;
	disk[1119] = 32'b00001100001001000000000000000000;
	disk[1120] = 32'b00101100000000010000000100110000;
	disk[1121] = 32'b00001100001001010000000000000000;
	disk[1122] = 32'b00110000000000010000000000000001;
	disk[1123] = 32'b00001100001000100000000000000000;
	disk[1124] = 32'b00001100101000110000000000000000;
	disk[1125] = 32'b00010000011000100000100000000000;
	disk[1126] = 32'b00001100001000100000000000000000;
	disk[1127] = 32'b00001100100000110000000000000000;
	disk[1128] = 32'b01011100011000100000010001101011;
	disk[1129] = 32'b00110000000000010000000000000000;
	disk[1130] = 32'b00110100000000010000000100101110;
	disk[1131] = 32'b00101100000000010000000100110000;
	disk[1132] = 32'b00001100001001000000000000000000;
	disk[1133] = 32'b00110000000000010000000000000001;
	disk[1134] = 32'b00001100001000100000000000000000;
	disk[1135] = 32'b00001100100000110000000000000000;
	disk[1136] = 32'b00010000011000100000100000000000;
	disk[1137] = 32'b00110100000000010000000100110000;
	disk[1138] = 32'b00111000000000000000010010011011;
	disk[1139] = 32'b00101100000000010000000100101110;
	disk[1140] = 32'b00001100001001000000000000000000;
	disk[1141] = 32'b00110000000000010000000000000000;
	disk[1142] = 32'b00001100001000100000000000000000;
	disk[1143] = 32'b00001100100000110000000000000000;
	disk[1144] = 32'b01011100011000100000010010000001;
	disk[1145] = 32'b00101100000000010000000100110000;
	disk[1146] = 32'b00001100001001000000000000000000;
	disk[1147] = 32'b00110000000000010000000000000001;
	disk[1148] = 32'b00001100001000100000000000000000;
	disk[1149] = 32'b00001100100000110000000000000000;
	disk[1150] = 32'b00010000011000100000100000000000;
	disk[1151] = 32'b00110100000000010000000100110100;
	disk[1152] = 32'b00111000000000000000010010001000;
	disk[1153] = 32'b00101100000000010000000100101110;
	disk[1154] = 32'b00001100001001000000000000000000;
	disk[1155] = 32'b00110000000000010000000000000001;
	disk[1156] = 32'b00001100001000100000000000000000;
	disk[1157] = 32'b00001100100000110000000000000000;
	disk[1158] = 32'b00010000011000100000100000000000;
	disk[1159] = 32'b00110100000000010000000100110100;
	disk[1160] = 32'b00101100000000010000000100110100;
	disk[1161] = 32'b00001100001001000000000000000000;
	disk[1162] = 32'b10100000000000010000000000000000;
	disk[1163] = 32'b00110100100000010000000011101101;
	disk[1164] = 32'b00001111110111101111111111111111;
	disk[1165] = 32'b00110111110111110000000000000000;
	disk[1166] = 32'b00101100000000010000000100110100;
	disk[1167] = 32'b00101100001000010000000011100011;
	disk[1168] = 32'b00001100001001000000000000000000;
	disk[1169] = 32'b00110000000000010000000000000001;
	disk[1170] = 32'b00001100001000100000000000000000;
	disk[1171] = 32'b00001100100000110000000000000000;
	disk[1172] = 32'b00010000011000100000100000000000;
	disk[1173] = 32'b00110100000000010000000101011011;
	disk[1174] = 32'b00101100000000010000000101011011;
	disk[1175] = 32'b00110100000000010000000100101010;
	disk[1176] = 32'b10000100000000000000001110000111;
	disk[1177] = 32'b00101111110111110000000000000000;
	disk[1178] = 32'b00001111110111100000000000000001;
	disk[1179] = 32'b00001111110111101111111111111111;
	disk[1180] = 32'b00110111110111110000000000000000;
	disk[1181] = 32'b00101100000000010000000100101110;
	disk[1182] = 32'b00101100001000010000000011100011;
	disk[1183] = 32'b00001100001001000000000000000000;
	disk[1184] = 32'b00110000000000010000000000000001;
	disk[1185] = 32'b00001100001000100000000000000000;
	disk[1186] = 32'b00001100100000110000000000000000;
	disk[1187] = 32'b00010000011000100000100000000000;
	disk[1188] = 32'b00110100000000010000000101011011;
	disk[1189] = 32'b00101100000000010000000101011011;
	disk[1190] = 32'b00110100000000010000000100101001;
	disk[1191] = 32'b10000100000000000000001101110001;
	disk[1192] = 32'b00101111110111110000000000000000;
	disk[1193] = 32'b00001111110111100000000000000001;
	disk[1194] = 32'b00001111110111101111111111111111;
	disk[1195] = 32'b00110111110111110000000000000000;
	disk[1196] = 32'b00101100000000010000000100101110;
	disk[1197] = 32'b00101100001000010000000011011001;
	disk[1198] = 32'b00110100000000010000000101011011;
	disk[1199] = 32'b00101100000000010000000101011011;
	disk[1200] = 32'b00110100000000010000000100100100;
	disk[1201] = 32'b10000100000000000000001100101000;
	disk[1202] = 32'b00101111110111110000000000000000;
	disk[1203] = 32'b00001111110111100000000000000001;
	disk[1204] = 32'b00101100000000010000000100101110;
	disk[1205] = 32'b00101100001000010000000011101101;
	disk[1206] = 32'b10100100001000000000000000000000;
	disk[1207] = 32'b00101100000000010000000100101110;
	disk[1208] = 32'b10000000001000000000000011101101;
	disk[1209] = 32'b00101100000000010000000100101110;
	disk[1210] = 32'b00101100001000010000000011100011;
	disk[1211] = 32'b00110100000000010000000100110101;
	disk[1212] = 32'b00101100000000010000000000000010;
	disk[1213] = 32'b00001100001001000000000000000000;
	disk[1214] = 32'b00110000000000010000000000000000;
	disk[1215] = 32'b00001100001000100000000000000000;
	disk[1216] = 32'b00001100100000110000000000000000;
	disk[1217] = 32'b01011100011000100000010011000011;
	disk[1218] = 32'b11000000000000000000000000000000;
	disk[1219] = 32'b00101100000000010000000000000010;
	disk[1220] = 32'b00001100001001000000000000000000;
	disk[1221] = 32'b00110000000000010000000000000011;
	disk[1222] = 32'b00001100001000100000000000000000;
	disk[1223] = 32'b00001100100000110000000000000000;
	disk[1224] = 32'b01011100011000100000010011001010;
	disk[1225] = 32'b11000000000000000000000000000000;
	disk[1226] = 32'b00101100000100110000000100110101;
	disk[1227] = 32'b10010100000100110000000000000000;
	disk[1228] = 32'b00101100000100110000000100110101;
	disk[1229] = 32'b10001100000100110000000000000000;
	disk[1230] = 32'b10101100000000000000000000000000;
	disk[1231] = 32'b00000000000000000000000000000000;
	disk[1232] = 32'b00110000000100110000000000000000;
	disk[1233] = 32'b10010100000100110000000000000000;
	disk[1234] = 32'b00110000000100110000000000000000;
	disk[1235] = 32'b10001100000100110000000000000000;
	disk[1236] = 32'b10101000000000000000100000000000;
	disk[1237] = 32'b00110100000000010000000000000010;
	disk[1238] = 32'b00101100000000010000000100101110;
	disk[1239] = 32'b00101100001000010000000011011001;
	disk[1240] = 32'b00110100000000010000000100110010;
	disk[1241] = 32'b00101100000000010000000100000100;
	disk[1242] = 32'b10011000001000000000000000000000;
	disk[1243] = 32'b10000000000000000000000100110010;
	disk[1244] = 32'b00101100000000010000000100000010;
	disk[1245] = 32'b10011000001000000000000000000000;
	disk[1246] = 32'b00101100000000010000000000000010;
	disk[1247] = 32'b00001100001001000000000000000000;
	disk[1248] = 32'b00110000000000010000000000000000;
	disk[1249] = 32'b00001100001000100000000000000000;
	disk[1250] = 32'b00001100100000110000000000000000;
	disk[1251] = 32'b01011100011000100000010011111110;
	disk[1252] = 32'b00110000000000010000000000000000;
	disk[1253] = 32'b00110100000000010000000100110011;
	disk[1254] = 32'b00110000000000010000000000000001;
	disk[1255] = 32'b00110100000000010000000100110001;
	disk[1256] = 32'b00101100000000010000000100101110;
	disk[1257] = 32'b00001100001001000000000000000000;
	disk[1258] = 32'b00101100000000010000000100110000;
	disk[1259] = 32'b00001100001001010000000000000000;
	disk[1260] = 32'b00110000000000010000000000000001;
	disk[1261] = 32'b00001100001000100000000000000000;
	disk[1262] = 32'b00001100101000110000000000000000;
	disk[1263] = 32'b00010000011000100000100000000000;
	disk[1264] = 32'b00001100001000100000000000000000;
	disk[1265] = 32'b00001100100000110000000000000000;
	disk[1266] = 32'b01011100011000100000010011110110;
	disk[1267] = 32'b00110000000000010000000000000000;
	disk[1268] = 32'b00110100000000010000000100101110;
	disk[1269] = 32'b00111000000000000000010011111101;
	disk[1270] = 32'b00101100000000010000000100101110;
	disk[1271] = 32'b00001100001001000000000000000000;
	disk[1272] = 32'b00110000000000010000000000000001;
	disk[1273] = 32'b00001100001000100000000000000000;
	disk[1274] = 32'b00001100100000110000000000000000;
	disk[1275] = 32'b00001000011000100000100000000000;
	disk[1276] = 32'b00110100000000010000000100101110;
	disk[1277] = 32'b00111000000000000000010100110000;
	disk[1278] = 32'b00101100000000010000000000000010;
	disk[1279] = 32'b00001100001001000000000000000000;
	disk[1280] = 32'b00110000000000010000000000000001;
	disk[1281] = 32'b00001100001000100000000000000000;
	disk[1282] = 32'b00001100100000110000000000000000;
	disk[1283] = 32'b01011100011000100000010100001110;
	disk[1284] = 32'b00110000000000010000000000000000;
	disk[1285] = 32'b00110100000000010000000100110011;
	disk[1286] = 32'b00110000000000010000000000000000;
	disk[1287] = 32'b00110100000000010000000100110001;
	disk[1288] = 32'b00001111110111101111111111111111;
	disk[1289] = 32'b00110111110111110000000000000000;
	disk[1290] = 32'b10000100000000000000001100011111;
	disk[1291] = 32'b00101111110111110000000000000000;
	disk[1292] = 32'b00001111110111100000000000000001;
	disk[1293] = 32'b00111000000000000000010100110000;
	disk[1294] = 32'b00101100000000010000000000000010;
	disk[1295] = 32'b00001100001001000000000000000000;
	disk[1296] = 32'b00110000000000010000000000000010;
	disk[1297] = 32'b00001100001000100000000000000000;
	disk[1298] = 32'b00001100100000110000000000000000;
	disk[1299] = 32'b01011100011000100000010100011110;
	disk[1300] = 32'b00110000000000010000000000000000;
	disk[1301] = 32'b00110100000000010000000100110011;
	disk[1302] = 32'b00110000000000010000000000000000;
	disk[1303] = 32'b00110100000000010000000100110001;
	disk[1304] = 32'b00001111110111101111111111111111;
	disk[1305] = 32'b00110111110111110000000000000000;
	disk[1306] = 32'b10000100000000000000001100100100;
	disk[1307] = 32'b00101111110111110000000000000000;
	disk[1308] = 32'b00001111110111100000000000000001;
	disk[1309] = 32'b00111000000000000000010100110000;
	disk[1310] = 32'b00101100000000010000000000000010;
	disk[1311] = 32'b00001100001001000000000000000000;
	disk[1312] = 32'b00110000000000010000000000000011;
	disk[1313] = 32'b00001100001000100000000000000000;
	disk[1314] = 32'b00001100100000110000000000000000;
	disk[1315] = 32'b01011100011000100000010100110000;
	disk[1316] = 32'b00110000000000010000000000000001;
	disk[1317] = 32'b00110100000000010000000100110011;
	disk[1318] = 32'b00110000000000010000000000000001;
	disk[1319] = 32'b00110100000000010000000100110001;
	disk[1320] = 32'b00101100000000010000000100110000;
	disk[1321] = 32'b00001100001001000000000000000000;
	disk[1322] = 32'b00110000000000010000000000000001;
	disk[1323] = 32'b00001100001000100000000000000000;
	disk[1324] = 32'b00001100100000110000000000000000;
	disk[1325] = 32'b01011100011000100000010100110000;
	disk[1326] = 32'b00110000000000010000000000000000;
	disk[1327] = 32'b00110100000000010000000100110000;
	disk[1328] = 32'b00111000000000000000010000001110;
	disk[1329] = 32'b00111111111000000000000000000000;
	disk[1330] = 32'b00110000000000010000000000001010;
	disk[1331] = 32'b00110100000000010000000100110110;
	disk[1332] = 32'b00101100000000010000000011111011;
	disk[1333] = 32'b10011000001000000000000000000000;
	disk[1334] = 32'b10000100000000000000000101011101;
	disk[1335] = 32'b00101100000000010000000100110110;
	disk[1336] = 32'b00001100001001000000000000000000;
	disk[1337] = 32'b00110000000000010000000000000000;
	disk[1338] = 32'b00001100001000100000000000000000;
	disk[1339] = 32'b00001100100000110000000000000000;
	disk[1340] = 32'b01100000011000100000010101100001;
	disk[1341] = 32'b00101100000000010000000011111011;
	disk[1342] = 32'b10011000001000000000000000000000;
	disk[1343] = 32'b01111100000000010000000000000000;
	disk[1344] = 32'b00110100000000010000000100110110;
	disk[1345] = 32'b00101100000000010000000100110110;
	disk[1346] = 32'b00001100001001000000000000000000;
	disk[1347] = 32'b00110000000000010000000000000001;
	disk[1348] = 32'b00001100001000100000000000000000;
	disk[1349] = 32'b00001100100000110000000000000000;
	disk[1350] = 32'b01011100011000100000010101001001;
	disk[1351] = 32'b10000100000000000000001001101110;
	disk[1352] = 32'b00111000000000000000010101100000;
	disk[1353] = 32'b00101100000000010000000100110110;
	disk[1354] = 32'b00001100001001000000000000000000;
	disk[1355] = 32'b00110000000000010000000000000010;
	disk[1356] = 32'b00001100001000100000000000000000;
	disk[1357] = 32'b00001100100000110000000000000000;
	disk[1358] = 32'b01011100011000100000010101010001;
	disk[1359] = 32'b10000100000000000000000110100101;
	disk[1360] = 32'b00111000000000000000010101100000;
	disk[1361] = 32'b00101100000000010000000100110110;
	disk[1362] = 32'b00001100001001000000000000000000;
	disk[1363] = 32'b00110000000000010000000000000011;
	disk[1364] = 32'b00001100001000100000000000000000;
	disk[1365] = 32'b00001100100000110000000000000000;
	disk[1366] = 32'b01011100011000100000010101011001;
	disk[1367] = 32'b10000100000000000000000111100000;
	disk[1368] = 32'b00111000000000000000010101100000;
	disk[1369] = 32'b00101100000000010000000100110110;
	disk[1370] = 32'b00001100001001000000000000000000;
	disk[1371] = 32'b00110000000000010000000000000100;
	disk[1372] = 32'b00001100001000100000000000000000;
	disk[1373] = 32'b00001100100000110000000000000000;
	disk[1374] = 32'b01011100011000100000010101100000;
	disk[1375] = 32'b10000100000000000000001111111001;
	disk[1376] = 32'b00111000000000000000010100110111;
	disk[1377] = 32'b00000100000000000000000000000000;


			// Program 1
			disk[1*(ADDR_WIDTH/TRACKS)+0] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+1] =  32'b00111000000000000000000000111001;
			disk[1*(ADDR_WIDTH/TRACKS)+2] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+3] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+4] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+5] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+6] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+7] =  32'b01110000011000100000000000001011;
			disk[1*(ADDR_WIDTH/TRACKS)+8] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+9] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+10] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+11] =  32'b00001111110111101111111111111110;
			disk[1*(ADDR_WIDTH/TRACKS)+12] =  32'b00110111110111110000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+13] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+14] =  32'b00110111110000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+15] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+16] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+17] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+18] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+19] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+20] =  32'b00010000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+21] =  32'b00110100000000010000000101011011;
			disk[1*(ADDR_WIDTH/TRACKS)+22] =  32'b00101100000000010000000101011011;
			disk[1*(ADDR_WIDTH/TRACKS)+23] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+24] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+25] =  32'b00101111110000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+26] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+27] =  32'b00101111110111110000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+28] =  32'b00001111110111100000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+29] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+30] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+31] =  32'b00001111110111101111111111111101;
			disk[1*(ADDR_WIDTH/TRACKS)+32] =  32'b00110111110111110000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+33] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+34] =  32'b00110111110000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+35] =  32'b00110111110001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+36] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+37] =  32'b00001100001001010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+38] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+39] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+40] =  32'b00001100101000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+41] =  32'b00010000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+42] =  32'b00110100000000010000000101011011;
			disk[1*(ADDR_WIDTH/TRACKS)+43] =  32'b00101100000000010000000101011011;
			disk[1*(ADDR_WIDTH/TRACKS)+44] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+45] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+46] =  32'b00101111110001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+47] =  32'b00101111110000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+48] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+49] =  32'b00101111110111110000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+50] =  32'b00001111110111100000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+51] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+52] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+53] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+54] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+55] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+56] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+57] =  32'b00110000000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+58] =  32'b00110100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+59] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+60] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+61] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+62] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+63] =  32'b00110100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+64] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+65] =  32'b10110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+66] =  32'b10101100000000000000000010000000;
			disk[1*(ADDR_WIDTH/TRACKS)+67] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+68] =  32'b10101100000000000000000011000000;
			disk[1*(ADDR_WIDTH/TRACKS)+69] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+70] =  32'b00000100000000000000000000000000;


			// Program 2
			
			disk[1*(ADDR_WIDTH/TRACKS)+71] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+72] =  32'b00111000000000000000000000110001;
			disk[1*(ADDR_WIDTH/TRACKS)+73] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+74] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+75] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+76] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+77] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+78] =  32'b01011100011000100000000000001011;
			disk[1*(ADDR_WIDTH/TRACKS)+79] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+80] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+81] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+82] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+83] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+84] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+85] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+86] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+87] =  32'b01011100011000100000000000010101;
			disk[1*(ADDR_WIDTH/TRACKS)+88] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+89] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+90] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+91] =  32'b00111000000000000000000000110001;
			disk[1*(ADDR_WIDTH/TRACKS)+92] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+93] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+94] =  32'b00001111110111101111111111111101;
			disk[1*(ADDR_WIDTH/TRACKS)+95] =  32'b00110111110111110000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+96] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+97] =  32'b00110111110000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+98] =  32'b00110111110001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+99] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+100] =  32'b00001100001001010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+101] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+102] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+103] =  32'b00001100101000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+104] =  32'b00010000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+105] =  32'b00110100000000010000000101011011;
			disk[1*(ADDR_WIDTH/TRACKS)+106] =  32'b00101100000000010000000101011011;
			disk[1*(ADDR_WIDTH/TRACKS)+107] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+108] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+109] =  32'b00101111110001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+110] =  32'b00101111110000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+111] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+112] =  32'b00101111110111110000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+113] =  32'b00001111110111100000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+114] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+115] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+116] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+117] =  32'b00011000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+118] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+119] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+120] =  32'b10101100000000000000000001000000;
			disk[1*(ADDR_WIDTH/TRACKS)+121] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+122] =  32'b10110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+123] =  32'b00110100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+124] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+125] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+126] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+127] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+128] =  32'b00110100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+129] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+130] =  32'b10110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+131] =  32'b10101100000000000000000010000000;
			disk[1*(ADDR_WIDTH/TRACKS)+132] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+133] =  32'b10101100000000000000000011000000;
			disk[1*(ADDR_WIDTH/TRACKS)+134] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+135] =  32'b00000100000000000000000000000000;

			// Program 3
			
			disk[1*(ADDR_WIDTH/TRACKS)+136] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+137] =  32'b00111000000000000000000000011110;
			disk[1*(ADDR_WIDTH/TRACKS)+138] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+139] =  32'b00110100000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+140] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+141] =  32'b00110100000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+142] =  32'b00101100000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+143] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+144] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+145] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+146] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+147] =  32'b01110000011000100000000000011011;
			disk[1*(ADDR_WIDTH/TRACKS)+148] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+149] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+150] =  32'b00101100000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+151] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+152] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+153] =  32'b00011000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+154] =  32'b00110100000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+155] =  32'b00101100000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+156] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+157] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+158] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+159] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+160] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+161] =  32'b00110100000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+162] =  32'b00111000000000000000000000000110;
			disk[1*(ADDR_WIDTH/TRACKS)+163] =  32'b00101100000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+164] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+165] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+166] =  32'b10101100000000000000000001000000;
			disk[1*(ADDR_WIDTH/TRACKS)+167] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+168] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+169] =  32'b10110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+170] =  32'b00110100000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+171] =  32'b10101100000000000000000001000000;
			disk[1*(ADDR_WIDTH/TRACKS)+172] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+173] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+174] =  32'b10110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+175] =  32'b00110100000000010000000000000110;
			disk[1*(ADDR_WIDTH/TRACKS)+176] =  32'b00101100000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+177] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+178] =  32'b00101100000000010000000000000110;
			disk[1*(ADDR_WIDTH/TRACKS)+179] =  32'b00110100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+180] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+181] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+182] =  32'b00110100000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+183] =  32'b00101100000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+184] =  32'b10110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+185] =  32'b10101100000000000000000010000000;
			disk[1*(ADDR_WIDTH/TRACKS)+186] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+187] =  32'b10101100000000000000000011000000;
			disk[1*(ADDR_WIDTH/TRACKS)+188] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+189] =  32'b00000100000000000000000000000000;

			
			
			// Program 4
			
			disk[1*(ADDR_WIDTH/TRACKS)+190] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+191] =  32'b00111000000000000000000000100110;
			disk[1*(ADDR_WIDTH/TRACKS)+192] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+193] =  32'b00110100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+194] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+195] =  32'b00110100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+196] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+197] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+198] =  32'b00101100000000010000000000010101;
			disk[1*(ADDR_WIDTH/TRACKS)+199] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+200] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+201] =  32'b01110000011000100000000000011110;
			disk[1*(ADDR_WIDTH/TRACKS)+202] =  32'b00101100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+203] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+204] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+205] =  32'b00101100000000100000000000010100;
			disk[1*(ADDR_WIDTH/TRACKS)+206] =  32'b00001000010000010000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+207] =  32'b00101100001000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+208] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+209] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+210] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+211] =  32'b00110100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+212] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+213] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+214] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+215] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+216] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+217] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+218] =  32'b00110100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+219] =  32'b00111000000000000000000000000110;
			disk[1*(ADDR_WIDTH/TRACKS)+220] =  32'b00101100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+221] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+222] =  32'b00101100000000010000000000010101;
			disk[1*(ADDR_WIDTH/TRACKS)+223] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+224] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+225] =  32'b00011100011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+226] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+227] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+228] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+229] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+230] =  32'b00110000000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+231] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+232] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+233] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+234] =  32'b00110000000000010000000000000111;
			disk[1*(ADDR_WIDTH/TRACKS)+235] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+236] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+237] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+238] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+239] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+240] =  32'b00110000000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+241] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+242] =  32'b00110000000000010000000000001100;
			disk[1*(ADDR_WIDTH/TRACKS)+243] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+244] =  32'b00110000000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+245] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+246] =  32'b00110000000000010000000000010010;
			disk[1*(ADDR_WIDTH/TRACKS)+247] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+248] =  32'b00110000000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+249] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+250] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+251] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+252] =  32'b00110000000000010000000000000110;
			disk[1*(ADDR_WIDTH/TRACKS)+253] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+254] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+255] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+256] =  32'b00110000000000010000000000000111;
			disk[1*(ADDR_WIDTH/TRACKS)+257] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+258] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+259] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+260] =  32'b00110000000000010000000000001000;
			disk[1*(ADDR_WIDTH/TRACKS)+261] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+262] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+263] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+264] =  32'b00110000000000010000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+265] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+266] =  32'b00110000000000010000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+267] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+268] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+269] =  32'b00110100000000010000000000010100;
			disk[1*(ADDR_WIDTH/TRACKS)+270] =  32'b00110000000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+271] =  32'b00110100000000010000000000010101;
			disk[1*(ADDR_WIDTH/TRACKS)+272] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+273] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+274] =  32'b00110100000000010000000000011000;
			disk[1*(ADDR_WIDTH/TRACKS)+275] =  32'b00101100000000010000000000011000;
			disk[1*(ADDR_WIDTH/TRACKS)+276] =  32'b10110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+277] =  32'b10101100000000000000000010000000;
			disk[1*(ADDR_WIDTH/TRACKS)+278] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+279] =  32'b10101100000000000000000011000000;
			disk[1*(ADDR_WIDTH/TRACKS)+280] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+281] =  32'b00000100000000000000000000000000;

			
			// Program 5
			
			disk[1*(ADDR_WIDTH/TRACKS)+282] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+283] =  32'b00111000000000000000000000101000;
			disk[1*(ADDR_WIDTH/TRACKS)+284] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+285] =  32'b00110100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+286] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+287] =  32'b00101100000000100000000000010100;
			disk[1*(ADDR_WIDTH/TRACKS)+288] =  32'b00001000010000010000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+289] =  32'b00101100001000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+290] =  32'b00110100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+291] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+292] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+293] =  32'b00101100000000010000000000010101;
			disk[1*(ADDR_WIDTH/TRACKS)+294] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+295] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+296] =  32'b01110000011000100000000000100101;
			disk[1*(ADDR_WIDTH/TRACKS)+297] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+298] =  32'b00101100000000100000000000010100;
			disk[1*(ADDR_WIDTH/TRACKS)+299] =  32'b00001000010000010000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+300] =  32'b00101100001000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+301] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+302] =  32'b00101100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+303] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+304] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+305] =  32'b01101100011000100000000000011101;
			disk[1*(ADDR_WIDTH/TRACKS)+306] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+307] =  32'b00101100000000100000000000010100;
			disk[1*(ADDR_WIDTH/TRACKS)+308] =  32'b00001000010000010000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+309] =  32'b00101100001000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+310] =  32'b00110100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+311] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+312] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+313] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+314] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+315] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+316] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+317] =  32'b00110100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+318] =  32'b00111000000000000000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+319] =  32'b00101100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+320] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+321] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+322] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+323] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+324] =  32'b00110000000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+325] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+326] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+327] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+328] =  32'b00110000000000010000000000000111;
			disk[1*(ADDR_WIDTH/TRACKS)+329] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+330] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+331] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+332] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+333] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+334] =  32'b00110000000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+335] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+336] =  32'b00110000000000010000000000001111;
			disk[1*(ADDR_WIDTH/TRACKS)+337] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+338] =  32'b00110000000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+339] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+340] =  32'b00110000000000010000000000010010;
			disk[1*(ADDR_WIDTH/TRACKS)+341] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+342] =  32'b00110000000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+343] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+344] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+345] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+346] =  32'b00110000000000010000000000000110;
			disk[1*(ADDR_WIDTH/TRACKS)+347] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+348] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+349] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+350] =  32'b00110000000000010000000000000111;
			disk[1*(ADDR_WIDTH/TRACKS)+351] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+352] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+353] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+354] =  32'b00110000000000010000000000001000;
			disk[1*(ADDR_WIDTH/TRACKS)+355] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+356] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+357] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+358] =  32'b00110000000000010000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+359] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+360] =  32'b00110000000000010000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+361] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+362] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+363] =  32'b00110100000000010000000000010100;
			disk[1*(ADDR_WIDTH/TRACKS)+364] =  32'b00110000000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+365] =  32'b00110100000000010000000000010101;
			disk[1*(ADDR_WIDTH/TRACKS)+366] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+367] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+368] =  32'b00110100000000010000000000011000;
			disk[1*(ADDR_WIDTH/TRACKS)+369] =  32'b00101100000000010000000000011000;
			disk[1*(ADDR_WIDTH/TRACKS)+370] =  32'b10110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+371] =  32'b10101100000000000000000010000000;
			disk[1*(ADDR_WIDTH/TRACKS)+372] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+373] =  32'b10101100000000000000000011000000;
			disk[1*(ADDR_WIDTH/TRACKS)+374] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+375] =  32'b00000100000000000000000000000000;


			// Program 6
			
			disk[1*(ADDR_WIDTH/TRACKS)+376] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+377] =  32'b00111000000000000000000000101000;
			disk[1*(ADDR_WIDTH/TRACKS)+378] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+379] =  32'b00110100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+380] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+381] =  32'b00101100000000100000000000010100;
			disk[1*(ADDR_WIDTH/TRACKS)+382] =  32'b00001000010000010000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+383] =  32'b00101100001000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+384] =  32'b00110100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+385] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+386] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+387] =  32'b00101100000000010000000000010101;
			disk[1*(ADDR_WIDTH/TRACKS)+388] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+389] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+390] =  32'b01110000011000100000000000100101;
			disk[1*(ADDR_WIDTH/TRACKS)+391] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+392] =  32'b00101100000000100000000000010100;
			disk[1*(ADDR_WIDTH/TRACKS)+393] =  32'b00001000010000010000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+394] =  32'b00101100001000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+395] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+396] =  32'b00101100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+397] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+398] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+399] =  32'b01110000011000100000000000011101;
			disk[1*(ADDR_WIDTH/TRACKS)+400] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+401] =  32'b00101100000000100000000000010100;
			disk[1*(ADDR_WIDTH/TRACKS)+402] =  32'b00001000010000010000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+403] =  32'b00101100001000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+404] =  32'b00110100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+405] =  32'b00101100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+406] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+407] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+408] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+409] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+410] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+411] =  32'b00110100000000010000000000010111;
			disk[1*(ADDR_WIDTH/TRACKS)+412] =  32'b00111000000000000000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+413] =  32'b00101100000000010000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+414] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+415] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+416] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+417] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+418] =  32'b00110000000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+419] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+420] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+421] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+422] =  32'b00110000000000010000000000000111;
			disk[1*(ADDR_WIDTH/TRACKS)+423] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+424] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+425] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+426] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+427] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+428] =  32'b00110000000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+429] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+430] =  32'b00110000000000010000000000001111;
			disk[1*(ADDR_WIDTH/TRACKS)+431] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+432] =  32'b00110000000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+433] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+434] =  32'b00110000000000010000000000010010;
			disk[1*(ADDR_WIDTH/TRACKS)+435] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+436] =  32'b00110000000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+437] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+438] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+439] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+440] =  32'b00110000000000010000000000000110;
			disk[1*(ADDR_WIDTH/TRACKS)+441] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+442] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+443] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+444] =  32'b00110000000000010000000000000111;
			disk[1*(ADDR_WIDTH/TRACKS)+445] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+446] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+447] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+448] =  32'b00110000000000010000000000001000;
			disk[1*(ADDR_WIDTH/TRACKS)+449] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+450] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+451] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+452] =  32'b00110000000000010000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+453] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+454] =  32'b00110000000000010000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+455] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+456] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+457] =  32'b00110100000000010000000000010100;
			disk[1*(ADDR_WIDTH/TRACKS)+458] =  32'b00110000000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+459] =  32'b00110100000000010000000000010101;
			disk[1*(ADDR_WIDTH/TRACKS)+460] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+461] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+462] =  32'b00110100000000010000000000011000;
			disk[1*(ADDR_WIDTH/TRACKS)+463] =  32'b00101100000000010000000000011000;
			disk[1*(ADDR_WIDTH/TRACKS)+464] =  32'b10110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+465] =  32'b10101100000000000000000010000000;
			disk[1*(ADDR_WIDTH/TRACKS)+466] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+467] =  32'b10101100000000000000000011000000;
			disk[1*(ADDR_WIDTH/TRACKS)+468] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+469] =  32'b00000100000000000000000000000000;


			// Program 7
			
			disk[1*(ADDR_WIDTH/TRACKS)+470] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+471] =  32'b00111000000000000000000000110011;
			disk[1*(ADDR_WIDTH/TRACKS)+472] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+473] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+474] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+475] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+476] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+477] =  32'b01011100011000100000000000001100;
			disk[1*(ADDR_WIDTH/TRACKS)+478] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+479] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+480] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+481] =  32'b00111000000000000000000000110011;
			disk[1*(ADDR_WIDTH/TRACKS)+482] =  32'b00001111110111101111111111111101;
			disk[1*(ADDR_WIDTH/TRACKS)+483] =  32'b00110111110111110000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+484] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+485] =  32'b00110111110000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+486] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+487] =  32'b00110111110000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+488] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+489] =  32'b00110100000000010000000101011011;
			disk[1*(ADDR_WIDTH/TRACKS)+490] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+491] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+492] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+493] =  32'b00001100001001010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+494] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+495] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+496] =  32'b00001100101000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+497] =  32'b00011100011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+498] =  32'b00001100001001010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+499] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+500] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+501] =  32'b00001100101000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+502] =  32'b00011000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+503] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+504] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+505] =  32'b00010000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+506] =  32'b00110100000000010000000101011010;
			disk[1*(ADDR_WIDTH/TRACKS)+507] =  32'b00101100000000010000000101011010;
			disk[1*(ADDR_WIDTH/TRACKS)+508] =  32'b00110100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+509] =  32'b00101100000000010000000101011011;
			disk[1*(ADDR_WIDTH/TRACKS)+510] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+511] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+512] =  32'b00101111110000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+513] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+514] =  32'b00101111110000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+515] =  32'b00110100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+516] =  32'b00101111110111110000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+517] =  32'b00001111110111100000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+518] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+519] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+520] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+521] =  32'b10101100000000000000000001000000;
			disk[1*(ADDR_WIDTH/TRACKS)+522] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+523] =  32'b10110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+524] =  32'b00110100000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+525] =  32'b10101100000000000000000001000000;
			disk[1*(ADDR_WIDTH/TRACKS)+526] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+527] =  32'b10110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+528] =  32'b00110100000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+529] =  32'b00101100000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+530] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+531] =  32'b00101100000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+532] =  32'b00110100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+533] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+534] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+535] =  32'b00110100000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+536] =  32'b00101100000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+537] =  32'b10110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+538] =  32'b10101100000000000000000010000000;
			disk[1*(ADDR_WIDTH/TRACKS)+539] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+540] =  32'b10101100000000000000000011000000;
			disk[1*(ADDR_WIDTH/TRACKS)+541] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+542] =  32'b00000100000000000000000000000000;


			// Program 8
			
			disk[1*(ADDR_WIDTH/TRACKS)+543] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+544] =  32'b00111000000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+545] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+546] =  32'b00110100000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+547] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+548] =  32'b00110100000000010000000000001011;
			disk[1*(ADDR_WIDTH/TRACKS)+549] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+550] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+551] =  32'b00110000000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+552] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+553] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+554] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+555] =  32'b00110000000000010000000000000111;
			disk[1*(ADDR_WIDTH/TRACKS)+556] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+557] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+558] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+559] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+560] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+561] =  32'b00110000000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+562] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+563] =  32'b00110000000000010000000000001111;
			disk[1*(ADDR_WIDTH/TRACKS)+564] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+565] =  32'b00110000000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+566] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+567] =  32'b00110000000000010000000000010010;
			disk[1*(ADDR_WIDTH/TRACKS)+568] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+569] =  32'b00110000000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+570] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+571] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+572] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+573] =  32'b00110000000000010000000000000110;
			disk[1*(ADDR_WIDTH/TRACKS)+574] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+575] =  32'b00110000000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+576] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+577] =  32'b00110000000000010000000000000111;
			disk[1*(ADDR_WIDTH/TRACKS)+578] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+579] =  32'b00110000000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+580] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+581] =  32'b00110000000000010000000000001000;
			disk[1*(ADDR_WIDTH/TRACKS)+582] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+583] =  32'b00110000000000010000000000011011;
			disk[1*(ADDR_WIDTH/TRACKS)+584] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+585] =  32'b00110000000000010000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+586] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+587] =  32'b00110000000000010000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+588] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+589] =  32'b00101100000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+590] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+591] =  32'b00110000000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+592] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+593] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+594] =  32'b01110000011000100000000001000100;
			disk[1*(ADDR_WIDTH/TRACKS)+595] =  32'b00101100000000010000000000001011;
			disk[1*(ADDR_WIDTH/TRACKS)+596] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+597] =  32'b00101100000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+598] =  32'b00101100001000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+599] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+600] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+601] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+602] =  32'b00110100000000010000000000001011;
			disk[1*(ADDR_WIDTH/TRACKS)+603] =  32'b00101100000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+604] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+605] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+606] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+607] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+608] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+609] =  32'b00110100000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+610] =  32'b00111000000000000000000000101110;
			disk[1*(ADDR_WIDTH/TRACKS)+611] =  32'b00101100000000010000000000001011;
			disk[1*(ADDR_WIDTH/TRACKS)+612] =  32'b10110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+613] =  32'b10101100000000000000000010000000;
			disk[1*(ADDR_WIDTH/TRACKS)+614] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+615] =  32'b10101100000000000000000011000000;
			disk[1*(ADDR_WIDTH/TRACKS)+616] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+617] =  32'b00000100000000000000000000000000;

			
			// Program 9
			
			disk[1*(ADDR_WIDTH/TRACKS)+618] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+619] =  32'b00111000000000000000000000100001;
			disk[1*(ADDR_WIDTH/TRACKS)+620] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+621] =  32'b00110100000000010000000000001101;
			disk[1*(ADDR_WIDTH/TRACKS)+622] =  32'b00101100000000010000000000001101;
			disk[1*(ADDR_WIDTH/TRACKS)+623] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+624] =  32'b00101100000000010000000000001011;
			disk[1*(ADDR_WIDTH/TRACKS)+625] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+626] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+627] =  32'b01110000011000100000000000011110;
			disk[1*(ADDR_WIDTH/TRACKS)+628] =  32'b00101100000000010000000000001101;
			disk[1*(ADDR_WIDTH/TRACKS)+629] =  32'b00101100000000100000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+630] =  32'b00001000010000010000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+631] =  32'b00101100001000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+632] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+633] =  32'b00101100000000010000000000001100;
			disk[1*(ADDR_WIDTH/TRACKS)+634] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+635] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+636] =  32'b01011100011000100000000000010110;
			disk[1*(ADDR_WIDTH/TRACKS)+637] =  32'b00101100000000010000000000001101;
			disk[1*(ADDR_WIDTH/TRACKS)+638] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+639] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+640] =  32'b00101100000000010000000000001101;
			disk[1*(ADDR_WIDTH/TRACKS)+641] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+642] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+643] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+644] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+645] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+646] =  32'b00110100000000010000000000001101;
			disk[1*(ADDR_WIDTH/TRACKS)+647] =  32'b00111000000000000000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+648] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+649] =  32'b00001100001111010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+650] =  32'b00111111111000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+651] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+652] =  32'b00110100000000010000000000001110;
			disk[1*(ADDR_WIDTH/TRACKS)+653] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+654] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+655] =  32'b00110000000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+656] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+657] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+658] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+659] =  32'b00110000000000010000000000000111;
			disk[1*(ADDR_WIDTH/TRACKS)+660] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+661] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+662] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+663] =  32'b00110000000000010000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+664] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+665] =  32'b00110000000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+666] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+667] =  32'b00110000000000010000000000001111;
			disk[1*(ADDR_WIDTH/TRACKS)+668] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+669] =  32'b00110000000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+670] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+671] =  32'b00110000000000010000000000010010;
			disk[1*(ADDR_WIDTH/TRACKS)+672] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+673] =  32'b00110000000000010000000000000101;
			disk[1*(ADDR_WIDTH/TRACKS)+674] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+675] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+676] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+677] =  32'b00110000000000010000000000000110;
			disk[1*(ADDR_WIDTH/TRACKS)+678] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+679] =  32'b00110000000000010000000000000011;
			disk[1*(ADDR_WIDTH/TRACKS)+680] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+681] =  32'b00110000000000010000000000000111;
			disk[1*(ADDR_WIDTH/TRACKS)+682] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+683] =  32'b00110000000000010000000000000100;
			disk[1*(ADDR_WIDTH/TRACKS)+684] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+685] =  32'b00110000000000010000000000001000;
			disk[1*(ADDR_WIDTH/TRACKS)+686] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+687] =  32'b00110000000000010000000000011011;
			disk[1*(ADDR_WIDTH/TRACKS)+688] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+689] =  32'b00110000000000010000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+690] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+691] =  32'b00110000000000010000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+692] =  32'b00110100100000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+693] =  32'b10101100000000000000000001000000;
			disk[1*(ADDR_WIDTH/TRACKS)+694] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+695] =  32'b10110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+696] =  32'b00110100000000010000000000001110;
			disk[1*(ADDR_WIDTH/TRACKS)+697] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+698] =  32'b00110100000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+699] =  32'b00110000000000010000000000001010;
			disk[1*(ADDR_WIDTH/TRACKS)+700] =  32'b00110100000000010000000000001011;
			disk[1*(ADDR_WIDTH/TRACKS)+701] =  32'b00101100000000010000000000001110;
			disk[1*(ADDR_WIDTH/TRACKS)+702] =  32'b00110100000000010000000000001100;
			disk[1*(ADDR_WIDTH/TRACKS)+703] =  32'b10000100000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+704] =  32'b00001111101000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+705] =  32'b00110100000000010000000000001110;
			disk[1*(ADDR_WIDTH/TRACKS)+706] =  32'b00101100000000010000000000001110;
			disk[1*(ADDR_WIDTH/TRACKS)+707] =  32'b10110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+708] =  32'b10101100000000000000000010000000;
			disk[1*(ADDR_WIDTH/TRACKS)+709] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+710] =  32'b10101100000000000000000011000000;
			disk[1*(ADDR_WIDTH/TRACKS)+711] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+712] =  32'b00000100000000000000000000000000;

			
			// Program 10

			disk[1*(ADDR_WIDTH/TRACKS)+713] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+714] =  32'b00111000000000000000000000000010;
			disk[1*(ADDR_WIDTH/TRACKS)+715] =  32'b00110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+716] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+717] =  32'b10101100000000000000000001000000;
			disk[1*(ADDR_WIDTH/TRACKS)+718] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+719] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+720] =  32'b10110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+721] =  32'b00110100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+722] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+723] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+724] =  32'b00110000000000010000000000001000;
			disk[1*(ADDR_WIDTH/TRACKS)+725] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+726] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+727] =  32'b01110000011000100000000000100011;
			disk[1*(ADDR_WIDTH/TRACKS)+728] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+729] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+730] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+731] =  32'b00001100001001010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+732] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+733] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+734] =  32'b00001100101000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+735] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+736] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+737] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+738] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+739] =  32'b00110100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+740] =  32'b00101100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+741] =  32'b00001100001001000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+742] =  32'b00110000000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+743] =  32'b00001100001000100000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+744] =  32'b00001100100000110000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+745] =  32'b00001000011000100000100000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+746] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+747] =  32'b00111000000000000000000000001001;
			disk[1*(ADDR_WIDTH/TRACKS)+748] =  32'b00101100000000010000000000000001;
			disk[1*(ADDR_WIDTH/TRACKS)+749] =  32'b10110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+750] =  32'b10101100000000000000000010000000;
			disk[1*(ADDR_WIDTH/TRACKS)+751] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+752] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+753] =  32'b10101100000000000000000001000000;
			disk[1*(ADDR_WIDTH/TRACKS)+754] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+755] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+756] =  32'b10110000000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+757] =  32'b00110100000000010000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+758] =  32'b10101100000000000000000011000000;
			disk[1*(ADDR_WIDTH/TRACKS)+759] =  32'b00000000000000000000000000000000;
			disk[1*(ADDR_WIDTH/TRACKS)+760] =  32'b00000100000000000000000000000000;


		end
	
	always @(posedge clock)
		begin
			if (hdFlag)
            begin
					disk[track*(ADDR_WIDTH/TRACKS) + trackPos] <= writeData;
            end
		end
		
		always@( posedge autoClock )
		begin
			readData <= disk[track*(ADDR_WIDTH/TRACKS) + trackPos];
		end
		

endmodule


