module InstructionMemory #(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=1000)
(adress, InstructionOut, clock, autoclock, rst);

	input [(DATA_WIDTH-1):0] adress;
	input clock, autoclock, rst;
	output reg [(DATA_WIDTH-1):0] InstructionOut;
	reg [(DATA_WIDTH-1):0] mem [ADDR_WIDTH-1:0];
	
	always @ (posedge clock)
		begin
			if( rst )
			begin
				mem[0] = 32'b00000000000000000000000000000000;
mem[1] = 32'b00111000000000000000001001011111;
mem[2] = 32'b00110000000000010000000000000000;
mem[3] = 32'b00110100000000010000000000010110;
mem[4] = 32'b00101100000000010000000000010110;
mem[5] = 32'b00001100001001000000000000000000;
mem[6] = 32'b00101100000000010000000000010101;
mem[7] = 32'b00001100001000100000000000000000;
mem[8] = 32'b00001100100000110000000000000000;
mem[9] = 32'b01110000011000100000000000011000;
mem[10] = 32'b00101100000000010000000000010110;
mem[11] = 32'b00101100000000100000000000010100;
mem[12] = 32'b00001000010000010000100000000000;
mem[13] = 32'b00001100001001000000000000000000;
mem[14] = 32'b01111100000000010000000000000000;
mem[15] = 32'b00110100100000010000000000000000;
mem[16] = 32'b00101100000000010000000000010110;
mem[17] = 32'b00001100001001000000000000000000;
mem[18] = 32'b00110000000000010000000000000001;
mem[19] = 32'b00001100001000100000000000000000;
mem[20] = 32'b00001100100000110000000000000000;
mem[21] = 32'b00001000011000100000100000000000;
mem[22] = 32'b00110100000000010000000000010110;
mem[23] = 32'b00111000000000000000000000000100;
mem[24] = 32'b00111111111000000000000000000000;
mem[25] = 32'b00110000000000010000000000000000;
mem[26] = 32'b00110100000000010000000000011001;
mem[27] = 32'b00101100000000010000000000011001;
mem[28] = 32'b00001100001001000000000000000000;
mem[29] = 32'b00101100000000010000000000011000;
mem[30] = 32'b00001100001000100000000000000000;
mem[31] = 32'b00001100100000110000000000000000;
mem[32] = 32'b01110000011000100000000000101111;
mem[33] = 32'b00101100000000010000000000011001;
mem[34] = 32'b00101100000000100000000000010111;
mem[35] = 32'b00001000010000010000100000000000;
mem[36] = 32'b00101100001000010000000000000000;
mem[37] = 32'b00110100000000010000000000011010;
mem[38] = 32'b10000000000000000000000000011010;
mem[39] = 32'b00101100000000010000000000011001;
mem[40] = 32'b00001100001001000000000000000000;
mem[41] = 32'b00110000000000010000000000000001;
mem[42] = 32'b00001100001000100000000000000000;
mem[43] = 32'b00001100100000110000000000000000;
mem[44] = 32'b00001000011000100000100000000000;
mem[45] = 32'b00110100000000010000000000011001;
mem[46] = 32'b00111000000000000000000000011011;
mem[47] = 32'b00111111111000000000000000000000;
mem[48] = 32'b00110000000000010000000000000001;
mem[49] = 32'b00110100000000010000000000011101;
mem[50] = 32'b00110000000000010000000000000000;
mem[51] = 32'b00110100000000010000000000011110;
mem[52] = 32'b00101100000000010000000000011110;
mem[53] = 32'b00001100001001000000000000000000;
mem[54] = 32'b00101100000000010000000000011100;
mem[55] = 32'b00001100001000100000000000000000;
mem[56] = 32'b00001100100000110000000000000000;
mem[57] = 32'b01110000011000100000000001001001;
mem[58] = 32'b00101100000000010000000000011011;
mem[59] = 32'b00001100001001000000000000000000;
mem[60] = 32'b00101100000000010000000000011101;
mem[61] = 32'b00001100001000100000000000000000;
mem[62] = 32'b00001100100000110000000000000000;
mem[63] = 32'b00011000011000100000100000000000;
mem[64] = 32'b00110100000000010000000000011101;
mem[65] = 32'b00101100000000010000000000011110;
mem[66] = 32'b00001100001001000000000000000000;
mem[67] = 32'b00110000000000010000000000000001;
mem[68] = 32'b00001100001000100000000000000000;
mem[69] = 32'b00001100100000110000000000000000;
mem[70] = 32'b00001000011000100000100000000000;
mem[71] = 32'b00110100000000010000000000011110;
mem[72] = 32'b00111000000000000000000000110100;
mem[73] = 32'b00101100000000010000000000011101;
mem[74] = 32'b00001100001111010000000000000000;
mem[75] = 32'b00111111111000000000000000000000;
mem[76] = 32'b00110000000000010000000000000000;
mem[77] = 32'b00110100000000010000000000100001;
mem[78] = 32'b00110000000000010000000000000000;
mem[79] = 32'b00110100000000010000000000100010;
mem[80] = 32'b00101100000000010000000000100010;
mem[81] = 32'b00001100001001000000000000000000;
mem[82] = 32'b00101100000000010000000000100000;
mem[83] = 32'b00001100001000100000000000000000;
mem[84] = 32'b00001100100000110000000000000000;
mem[85] = 32'b01110000011000100000000001101000;
mem[86] = 32'b00101100000000010000000000100001;
mem[87] = 32'b00001100001001000000000000000000;
mem[88] = 32'b00101100000000010000000000100010;
mem[89] = 32'b00101100000000100000000000011111;
mem[90] = 32'b00001000010000010000100000000000;
mem[91] = 32'b00101100001000010000000000000000;
mem[92] = 32'b00001100001000100000000000000000;
mem[93] = 32'b00001100100000110000000000000000;
mem[94] = 32'b00001000011000100000100000000000;
mem[95] = 32'b00110100000000010000000000100001;
mem[96] = 32'b00101100000000010000000000100010;
mem[97] = 32'b00001100001001000000000000000000;
mem[98] = 32'b00110000000000010000000000000001;
mem[99] = 32'b00001100001000100000000000000000;
mem[100] = 32'b00001100100000110000000000000000;
mem[101] = 32'b00001000011000100000100000000000;
mem[102] = 32'b00110100000000010000000000100010;
mem[103] = 32'b00111000000000000000000001010000;
mem[104] = 32'b00101100000000010000000000100001;
mem[105] = 32'b00001100001001000000000000000000;
mem[106] = 32'b00101100000000010000000000100000;
mem[107] = 32'b00001100001000100000000000000000;
mem[108] = 32'b00001100100000110000000000000000;
mem[109] = 32'b00011100011000100000100000000000;
mem[110] = 32'b00001100001111010000000000000000;
mem[111] = 32'b00111111111000000000000000000000;
mem[112] = 32'b00101100000000010000000000100100;
mem[113] = 32'b00001100001001000000000000000000;
mem[114] = 32'b00101100000000010000000000100101;
mem[115] = 32'b00001100001000100000000000000000;
mem[116] = 32'b00001100100000110000000000000000;
mem[117] = 32'b00001000011000100000100000000000;
mem[118] = 32'b00001100001001000000000000000000;
mem[119] = 32'b00110000000000010000000000000010;
mem[120] = 32'b00001100001000100000000000000000;
mem[121] = 32'b00001100100000110000000000000000;
mem[122] = 32'b00011100011000100000100000000000;
mem[123] = 32'b00110100000000010000000000100111;
mem[124] = 32'b00101100000000010000000000100101;
mem[125] = 32'b00001100001001000000000000000000;
mem[126] = 32'b00101100000000010000000000100100;
mem[127] = 32'b00001100001000100000000000000000;
mem[128] = 32'b00001100100000110000000000000000;
mem[129] = 32'b01110000011000100000000100001011;
mem[130] = 32'b00101100000000010000000000100111;
mem[131] = 32'b00001100001001000000000000000000;
mem[132] = 32'b00110000000000010000000000000001;
mem[133] = 32'b00001100001000100000000000000000;
mem[134] = 32'b00001100100000110000000000000000;
mem[135] = 32'b00010000011000100000100000000000;
mem[136] = 32'b00101100000000100000000000100011;
mem[137] = 32'b00001000010000010000100000000000;
mem[138] = 32'b00101100001000010000000000000000;
mem[139] = 32'b00001100001001000000000000000000;
mem[140] = 32'b00101100000000010000000000100110;
mem[141] = 32'b00001100001000100000000000000000;
mem[142] = 32'b00001100100000110000000000000000;
mem[143] = 32'b01011100011000100000000010010011;
mem[144] = 32'b00101100000000010000000000100111;
mem[145] = 32'b00001100001111010000000000000000;
mem[146] = 32'b00111111111000000000000000000000;
mem[147] = 32'b00101100000000010000000000100110;
mem[148] = 32'b00001100001001000000000000000000;
mem[149] = 32'b00101100000000010000000000100111;
mem[150] = 32'b00001100001001010000000000000000;
mem[151] = 32'b00110000000000010000000000000001;
mem[152] = 32'b00001100001000100000000000000000;
mem[153] = 32'b00001100101000110000000000000000;
mem[154] = 32'b00010000011000100000100000000000;
mem[155] = 32'b00101100000000100000000000100011;
mem[156] = 32'b00001000010000010000100000000000;
mem[157] = 32'b00101100001000010000000000000000;
mem[158] = 32'b00001100001000100000000000000000;
mem[159] = 32'b00001100100000110000000000000000;
mem[160] = 32'b01101100011000100000000011001111;
mem[161] = 32'b00001111110111101111111111111011;
mem[162] = 32'b00110111110111110000000000000100;
mem[163] = 32'b00101100000000010000000000100110;
mem[164] = 32'b00110111110000010000000000000011;
mem[165] = 32'b00101100000000010000000000100011;
mem[166] = 32'b00110111110000010000000000000010;
mem[167] = 32'b00101100000000010000000000100100;
mem[168] = 32'b00110111110000010000000000000001;
mem[169] = 32'b00101100000000010000000000100101;
mem[170] = 32'b00110111110000010000000000000000;
mem[171] = 32'b00101100000000010000000000100011;
mem[172] = 32'b00110100000000010000001111111110;
mem[173] = 32'b00101100000000010000000000100111;
mem[174] = 32'b00001100001001000000000000000000;
mem[175] = 32'b00110000000000010000000000000001;
mem[176] = 32'b00001100001000100000000000000000;
mem[177] = 32'b00001100100000110000000000000000;
mem[178] = 32'b00001000011000100000100000000000;
mem[179] = 32'b00110100000000010000001111111101;
mem[180] = 32'b00101100000000010000000000100101;
mem[181] = 32'b00110100000000010000001111111100;
mem[182] = 32'b00101100000000010000000000100110;
mem[183] = 32'b00110100000000010000001111111011;
mem[184] = 32'b00101100000000010000001111111011;
mem[185] = 32'b00110100000000010000000000100110;
mem[186] = 32'b00101100000000010000001111111100;
mem[187] = 32'b00110100000000010000000000100101;
mem[188] = 32'b00101100000000010000001111111101;
mem[189] = 32'b00110100000000010000000000100100;
mem[190] = 32'b00101100000000010000001111111110;
mem[191] = 32'b00110100000000010000000000100011;
mem[192] = 32'b10000100000000000000000001110000;
mem[193] = 32'b00101111110000010000000000000011;
mem[194] = 32'b00110100000000010000000000100110;
mem[195] = 32'b00101111110000010000000000000010;
mem[196] = 32'b00110100000000010000000000100011;
mem[197] = 32'b00101111110000010000000000000001;
mem[198] = 32'b00110100000000010000000000100100;
mem[199] = 32'b00101111110000010000000000000000;
mem[200] = 32'b00110100000000010000000000100101;
mem[201] = 32'b00101111110111110000000000000100;
mem[202] = 32'b00001111110111100000000000000101;
mem[203] = 32'b00001111101000010000000000000000;
mem[204] = 32'b00001100001111010000000000000000;
mem[205] = 32'b00111111111000000000000000000000;
mem[206] = 32'b00111000000000000000000100001001;
mem[207] = 32'b00101100000000010000000000100110;
mem[208] = 32'b00001100001001000000000000000000;
mem[209] = 32'b00101100000000010000000000100111;
mem[210] = 32'b00001100001001010000000000000000;
mem[211] = 32'b00110000000000010000000000000001;
mem[212] = 32'b00001100001000100000000000000000;
mem[213] = 32'b00001100101000110000000000000000;
mem[214] = 32'b00010000011000100000100000000000;
mem[215] = 32'b00101100000000100000000000100011;
mem[216] = 32'b00001000010000010000100000000000;
mem[217] = 32'b00101100001000010000000000000000;
mem[218] = 32'b00001100001000100000000000000000;
mem[219] = 32'b00001100100000110000000000000000;
mem[220] = 32'b01110000011000100000000100001010;
mem[221] = 32'b00001111110111101111111111111011;
mem[222] = 32'b00110111110111110000000000000100;
mem[223] = 32'b00101100000000010000000000100110;
mem[224] = 32'b00110111110000010000000000000011;
mem[225] = 32'b00101100000000010000000000100011;
mem[226] = 32'b00110111110000010000000000000010;
mem[227] = 32'b00101100000000010000000000100100;
mem[228] = 32'b00110111110000010000000000000001;
mem[229] = 32'b00101100000000010000000000100101;
mem[230] = 32'b00110111110000010000000000000000;
mem[231] = 32'b00101100000000010000000000100011;
mem[232] = 32'b00110100000000010000001111111110;
mem[233] = 32'b00101100000000010000000000100100;
mem[234] = 32'b00110100000000010000001111111101;
mem[235] = 32'b00101100000000010000000000100111;
mem[236] = 32'b00001100001001000000000000000000;
mem[237] = 32'b00110000000000010000000000000001;
mem[238] = 32'b00001100001000100000000000000000;
mem[239] = 32'b00001100100000110000000000000000;
mem[240] = 32'b00010000011000100000100000000000;
mem[241] = 32'b00110100000000010000001111111100;
mem[242] = 32'b00101100000000010000000000100110;
mem[243] = 32'b00110100000000010000001111111011;
mem[244] = 32'b00101100000000010000001111111011;
mem[245] = 32'b00110100000000010000000000100110;
mem[246] = 32'b00101100000000010000001111111100;
mem[247] = 32'b00110100000000010000000000100101;
mem[248] = 32'b00101100000000010000001111111101;
mem[249] = 32'b00110100000000010000000000100100;
mem[250] = 32'b00101100000000010000001111111110;
mem[251] = 32'b00110100000000010000000000100011;
mem[252] = 32'b10000100000000000000000001110000;
mem[253] = 32'b00101111110000010000000000000011;
mem[254] = 32'b00110100000000010000000000100110;
mem[255] = 32'b00101111110000010000000000000010;
mem[256] = 32'b00110100000000010000000000100011;
mem[257] = 32'b00101111110000010000000000000001;
mem[258] = 32'b00110100000000010000000000100100;
mem[259] = 32'b00101111110000010000000000000000;
mem[260] = 32'b00110100000000010000000000100101;
mem[261] = 32'b00101111110111110000000000000100;
mem[262] = 32'b00001111110111100000000000000101;
mem[263] = 32'b00001111101000010000000000000000;
mem[264] = 32'b00001100001111010000000000000000;
mem[265] = 32'b00111111111000000000000000000000;
mem[266] = 32'b00111000000000000000000100001101;
mem[267] = 32'b00110000000000010000000000000000;
mem[268] = 32'b00001100001111010000000000000000;
mem[269] = 32'b00111111111000000000000000000000;
mem[270] = 32'b00110000000000010000000000000000;
mem[271] = 32'b00110100000000010000000000101011;
mem[272] = 32'b00101100000000010000000000101011;
mem[273] = 32'b00101100000000100000000000101000;
mem[274] = 32'b00001000010000010000100000000000;
mem[275] = 32'b00101100001000010000000000000000;
mem[276] = 32'b00110100000000010000000000101010;
mem[277] = 32'b00101100000000010000000000101011;
mem[278] = 32'b00001100001001000000000000000000;
mem[279] = 32'b00101100000000010000000000101001;
mem[280] = 32'b00001100001000100000000000000000;
mem[281] = 32'b00001100100000110000000000000000;
mem[282] = 32'b01110000011000100000000100110001;
mem[283] = 32'b00101100000000010000000000101011;
mem[284] = 32'b00101100000000100000000000101000;
mem[285] = 32'b00001000010000010000100000000000;
mem[286] = 32'b00101100001000010000000000000000;
mem[287] = 32'b00001100001001000000000000000000;
mem[288] = 32'b00101100000000010000000000101010;
mem[289] = 32'b00001100001000100000000000000000;
mem[290] = 32'b00001100100000110000000000000000;
mem[291] = 32'b01101100011000100000000100101001;
mem[292] = 32'b00101100000000010000000000101011;
mem[293] = 32'b00101100000000100000000000101000;
mem[294] = 32'b00001000010000010000100000000000;
mem[295] = 32'b00101100001000010000000000000000;
mem[296] = 32'b00110100000000010000000000101010;
mem[297] = 32'b00101100000000010000000000101011;
mem[298] = 32'b00001100001001000000000000000000;
mem[299] = 32'b00110000000000010000000000000001;
mem[300] = 32'b00001100001000100000000000000000;
mem[301] = 32'b00001100100000110000000000000000;
mem[302] = 32'b00001000011000100000100000000000;
mem[303] = 32'b00110100000000010000000000101011;
mem[304] = 32'b00111000000000000000000100010101;
mem[305] = 32'b00101100000000010000000000101010;
mem[306] = 32'b00001100001111010000000000000000;
mem[307] = 32'b00111111111000000000000000000000;
mem[308] = 32'b00110000000000010000000000000000;
mem[309] = 32'b00110100000000010000000000101111;
mem[310] = 32'b00101100000000010000000000101111;
mem[311] = 32'b00101100000000100000000000101100;
mem[312] = 32'b00001000010000010000100000000000;
mem[313] = 32'b00101100001000010000000000000000;
mem[314] = 32'b00110100000000010000000000101110;
mem[315] = 32'b00101100000000010000000000101111;
mem[316] = 32'b00001100001001000000000000000000;
mem[317] = 32'b00101100000000010000000000101101;
mem[318] = 32'b00001100001000100000000000000000;
mem[319] = 32'b00001100100000110000000000000000;
mem[320] = 32'b01110000011000100000000101010111;
mem[321] = 32'b00101100000000010000000000101111;
mem[322] = 32'b00101100000000100000000000101100;
mem[323] = 32'b00001000010000010000100000000000;
mem[324] = 32'b00101100001000010000000000000000;
mem[325] = 32'b00001100001001000000000000000000;
mem[326] = 32'b00101100000000010000000000101110;
mem[327] = 32'b00001100001000100000000000000000;
mem[328] = 32'b00001100100000110000000000000000;
mem[329] = 32'b01110000011000100000000101001111;
mem[330] = 32'b00101100000000010000000000101111;
mem[331] = 32'b00101100000000100000000000101100;
mem[332] = 32'b00001000010000010000100000000000;
mem[333] = 32'b00101100001000010000000000000000;
mem[334] = 32'b00110100000000010000000000101110;
mem[335] = 32'b00101100000000010000000000101111;
mem[336] = 32'b00001100001001000000000000000000;
mem[337] = 32'b00110000000000010000000000000001;
mem[338] = 32'b00001100001000100000000000000000;
mem[339] = 32'b00001100100000110000000000000000;
mem[340] = 32'b00001000011000100000100000000000;
mem[341] = 32'b00110100000000010000000000101111;
mem[342] = 32'b00111000000000000000000100111011;
mem[343] = 32'b00101100000000010000000000101110;
mem[344] = 32'b00001100001111010000000000000000;
mem[345] = 32'b00111111111000000000000000000000;
mem[346] = 32'b00101100000000010000000000110000;
mem[347] = 32'b00001100001001000000000000000000;
mem[348] = 32'b00110000000000010000000000000010;
mem[349] = 32'b00001100001000100000000000000000;
mem[350] = 32'b00001100100000110000000000000000;
mem[351] = 32'b01110000011000100000000101100011;
mem[352] = 32'b00110000000000010000000000000001;
mem[353] = 32'b00001100001111010000000000000000;
mem[354] = 32'b00111111111000000000000000000000;
mem[355] = 32'b00001111110111101111111111111110;
mem[356] = 32'b00110111110111110000000000000001;
mem[357] = 32'b00101100000000010000000000110000;
mem[358] = 32'b00110111110000010000000000000000;
mem[359] = 32'b00101100000000010000000000110000;
mem[360] = 32'b00001100001001000000000000000000;
mem[361] = 32'b00110000000000010000000000000001;
mem[362] = 32'b00001100001000100000000000000000;
mem[363] = 32'b00001100100000110000000000000000;
mem[364] = 32'b00010000011000100000100000000000;
mem[365] = 32'b00110100000000010000001111111110;
mem[366] = 32'b00101100000000010000001111111110;
mem[367] = 32'b00110100000000010000000000110000;
mem[368] = 32'b10000100000000000000000101011010;
mem[369] = 32'b00101111110000010000000000000000;
mem[370] = 32'b00110100000000010000000000110000;
mem[371] = 32'b00101111110111110000000000000001;
mem[372] = 32'b00001111110111100000000000000010;
mem[373] = 32'b00001111101000010000000000000000;
mem[374] = 32'b00001100001001000000000000000000;
mem[375] = 32'b00001111110111101111111111111101;
mem[376] = 32'b00110111110111110000000000000010;
mem[377] = 32'b00101100000000010000000000110000;
mem[378] = 32'b00110111110000010000000000000001;
mem[379] = 32'b00110111110001000000000000000000;
mem[380] = 32'b00101100000000010000000000110000;
mem[381] = 32'b00001100001001010000000000000000;
mem[382] = 32'b00110000000000010000000000000010;
mem[383] = 32'b00001100001000100000000000000000;
mem[384] = 32'b00001100101000110000000000000000;
mem[385] = 32'b00010000011000100000100000000000;
mem[386] = 32'b00110100000000010000001111111110;
mem[387] = 32'b00101100000000010000001111111110;
mem[388] = 32'b00110100000000010000000000110000;
mem[389] = 32'b10000100000000000000000101011010;
mem[390] = 32'b00101111110001000000000000000000;
mem[391] = 32'b00101111110000010000000000000001;
mem[392] = 32'b00110100000000010000000000110000;
mem[393] = 32'b00101111110111110000000000000010;
mem[394] = 32'b00001111110111100000000000000011;
mem[395] = 32'b00001111101000010000000000000000;
mem[396] = 32'b00001100001000100000000000000000;
mem[397] = 32'b00001100100000110000000000000000;
mem[398] = 32'b00001000011000100000100000000000;
mem[399] = 32'b00001100001111010000000000000000;
mem[400] = 32'b00111111111000000000000000000000;
mem[401] = 32'b00101100000000010000000000110001;
mem[402] = 32'b00001100001001000000000000000000;
mem[403] = 32'b00110000000000010000000000000000;
mem[404] = 32'b00001100001000100000000000000000;
mem[405] = 32'b00001100100000110000000000000000;
mem[406] = 32'b01011100011000100000000110011010;
mem[407] = 32'b00110000000000010000000000000001;
mem[408] = 32'b00001100001111010000000000000000;
mem[409] = 32'b00111111111000000000000000000000;
mem[410] = 32'b00101100000000010000000000110001;
mem[411] = 32'b00001100001001000000000000000000;
mem[412] = 32'b00110000000000010000000000000001;
mem[413] = 32'b00001100001000100000000000000000;
mem[414] = 32'b00001100100000110000000000000000;
mem[415] = 32'b01011100011000100000000110100100;
mem[416] = 32'b00110000000000010000000000000001;
mem[417] = 32'b00001100001111010000000000000000;
mem[418] = 32'b00111111111000000000000000000000;
mem[419] = 32'b00111000000000000000000110111111;
mem[420] = 32'b00101100000000010000000000110001;
mem[421] = 32'b00001100001001000000000000000000;
mem[422] = 32'b00001111110111101111111111111101;
mem[423] = 32'b00110111110111110000000000000010;
mem[424] = 32'b00101100000000010000000000110001;
mem[425] = 32'b00110111110000010000000000000001;
mem[426] = 32'b00110111110001000000000000000000;
mem[427] = 32'b00101100000000010000000000110001;
mem[428] = 32'b00001100001001010000000000000000;
mem[429] = 32'b00110000000000010000000000000001;
mem[430] = 32'b00001100001000100000000000000000;
mem[431] = 32'b00001100101000110000000000000000;
mem[432] = 32'b00010000011000100000100000000000;
mem[433] = 32'b00110100000000010000001111111110;
mem[434] = 32'b00101100000000010000001111111110;
mem[435] = 32'b00110100000000010000000000110001;
mem[436] = 32'b10000100000000000000000110010001;
mem[437] = 32'b00101111110001000000000000000000;
mem[438] = 32'b00101111110000010000000000000001;
mem[439] = 32'b00110100000000010000000000110001;
mem[440] = 32'b00101111110111110000000000000010;
mem[441] = 32'b00001111110111100000000000000011;
mem[442] = 32'b00001111101000010000000000000000;
mem[443] = 32'b00001100001000100000000000000000;
mem[444] = 32'b00001100100000110000000000000000;
mem[445] = 32'b00011000011000100000100000000000;
mem[446] = 32'b00001100001111010000000000000000;
mem[447] = 32'b00111111111000000000000000000000;
mem[448] = 32'b10000000000000000000000000110010;
mem[449] = 32'b10000000000000000000000000110011;
mem[450] = 32'b00101100000000010000000000110011;
mem[451] = 32'b00001100001001000000000000000000;
mem[452] = 32'b00110000000000010000000000000000;
mem[453] = 32'b00001100001000100000000000000000;
mem[454] = 32'b00001100100000110000000000000000;
mem[455] = 32'b01011100011000100000000111001100;
mem[456] = 32'b00101100000000010000000000110010;
mem[457] = 32'b00001100001111010000000000000000;
mem[458] = 32'b00111111111000000000000000000000;
mem[459] = 32'b00111000000000000000000111110010;
mem[460] = 32'b00001111110111101111111111111101;
mem[461] = 32'b00110111110111110000000000000010;
mem[462] = 32'b00101100000000010000000000110010;
mem[463] = 32'b00110111110000010000000000000001;
mem[464] = 32'b00101100000000010000000000110011;
mem[465] = 32'b00110111110000010000000000000000;
mem[466] = 32'b00101100000000010000000000110011;
mem[467] = 32'b00110100000000010000001111111110;
mem[468] = 32'b00101100000000010000000000110010;
mem[469] = 32'b00001100001001000000000000000000;
mem[470] = 32'b00101100000000010000000000110010;
mem[471] = 32'b00001100001001010000000000000000;
mem[472] = 32'b00101100000000010000000000110011;
mem[473] = 32'b00001100001000100000000000000000;
mem[474] = 32'b00001100101000110000000000000000;
mem[475] = 32'b00011100011000100000100000000000;
mem[476] = 32'b00001100001001010000000000000000;
mem[477] = 32'b00101100000000010000000000110011;
mem[478] = 32'b00001100001000100000000000000000;
mem[479] = 32'b00001100101000110000000000000000;
mem[480] = 32'b00011000011000100000100000000000;
mem[481] = 32'b00001100001000100000000000000000;
mem[482] = 32'b00001100100000110000000000000000;
mem[483] = 32'b00010000011000100000100000000000;
mem[484] = 32'b00110100000000010000001111111101;
mem[485] = 32'b00101100000000010000001111111101;
mem[486] = 32'b00110100000000010000000000110011;
mem[487] = 32'b00101100000000010000001111111110;
mem[488] = 32'b00110100000000010000000000110010;
mem[489] = 32'b10000100000000000000000111000000;
mem[490] = 32'b00101111110000010000000000000001;
mem[491] = 32'b00110100000000010000000000110010;
mem[492] = 32'b00101111110000010000000000000000;
mem[493] = 32'b00110100000000010000000000110011;
mem[494] = 32'b00101111110111110000000000000010;
mem[495] = 32'b00001111110111100000000000000011;
mem[496] = 32'b00001111101000010000000000000000;
mem[497] = 32'b00001100001111010000000000000000;
mem[498] = 32'b00111111111000000000000000000000;
mem[499] = 32'b00101100000000010000000000110101;
mem[500] = 32'b00110100000000010000000000111001;
mem[501] = 32'b00101100000000010000000000110101;
mem[502] = 32'b00101100000000100000000000110100;
mem[503] = 32'b00001000010000010000100000000000;
mem[504] = 32'b00101100001000010000000000000000;
mem[505] = 32'b00110100000000010000000000111000;
mem[506] = 32'b00101100000000010000000000110101;
mem[507] = 32'b00001100001001000000000000000000;
mem[508] = 32'b00110000000000010000000000000001;
mem[509] = 32'b00001100001000100000000000000000;
mem[510] = 32'b00001100100000110000000000000000;
mem[511] = 32'b00001000011000100000100000000000;
mem[512] = 32'b00110100000000010000000000110111;
mem[513] = 32'b00101100000000010000000000110111;
mem[514] = 32'b00001100001001000000000000000000;
mem[515] = 32'b00101100000000010000000000110110;
mem[516] = 32'b00001100001000100000000000000000;
mem[517] = 32'b00001100100000110000000000000000;
mem[518] = 32'b01110000011000100000001000011111;
mem[519] = 32'b00101100000000010000000000110111;
mem[520] = 32'b00101100000000100000000000110100;
mem[521] = 32'b00001000010000010000100000000000;
mem[522] = 32'b00101100001000010000000000000000;
mem[523] = 32'b00001100001001000000000000000000;
mem[524] = 32'b00101100000000010000000000111000;
mem[525] = 32'b00001100001000100000000000000000;
mem[526] = 32'b00001100100000110000000000000000;
mem[527] = 32'b01110000011000100000001000010111;
mem[528] = 32'b00101100000000010000000000110111;
mem[529] = 32'b00101100000000100000000000110100;
mem[530] = 32'b00001000010000010000100000000000;
mem[531] = 32'b00101100001000010000000000000000;
mem[532] = 32'b00110100000000010000000000111000;
mem[533] = 32'b00101100000000010000000000110111;
mem[534] = 32'b00110100000000010000000000111001;
mem[535] = 32'b00101100000000010000000000110111;
mem[536] = 32'b00001100001001000000000000000000;
mem[537] = 32'b00110000000000010000000000000001;
mem[538] = 32'b00001100001000100000000000000000;
mem[539] = 32'b00001100100000110000000000000000;
mem[540] = 32'b00001000011000100000100000000000;
mem[541] = 32'b00110100000000010000000000110111;
mem[542] = 32'b00111000000000000000001000000001;
mem[543] = 32'b00101100000000010000000000111001;
mem[544] = 32'b00001100001111010000000000000000;
mem[545] = 32'b00111111111000000000000000000000;
mem[546] = 32'b00101100000000010000000000111011;
mem[547] = 32'b00110100000000010000000000111101;
mem[548] = 32'b00101100000000010000000000111101;
mem[549] = 32'b00001100001001000000000000000000;
mem[550] = 32'b00101100000000010000000000111100;
mem[551] = 32'b00001100001001010000000000000000;
mem[552] = 32'b00110000000000010000000000000001;
mem[553] = 32'b00001100001000100000000000000000;
mem[554] = 32'b00001100101000110000000000000000;
mem[555] = 32'b00010000011000100000100000000000;
mem[556] = 32'b00001100001000100000000000000000;
mem[557] = 32'b00001100100000110000000000000000;
mem[558] = 32'b01110000011000100000001001011110;
mem[559] = 32'b00001111110111101111111111111111;
mem[560] = 32'b00110111110111110000000000000000;
mem[561] = 32'b00101100000000010000000000111010;
mem[562] = 32'b00110100000000010000001111111110;
mem[563] = 32'b00101100000000010000000000111101;
mem[564] = 32'b00110100000000010000001111111101;
mem[565] = 32'b00101100000000010000000000111100;
mem[566] = 32'b00110100000000010000001111111100;
mem[567] = 32'b00101100000000010000001111111100;
mem[568] = 32'b00110100000000010000000000110110;
mem[569] = 32'b00101100000000010000001111111101;
mem[570] = 32'b00110100000000010000000000110101;
mem[571] = 32'b00101100000000010000001111111110;
mem[572] = 32'b00110100000000010000000000110100;
mem[573] = 32'b10000100000000000000000111110011;
mem[574] = 32'b00101111110111110000000000000000;
mem[575] = 32'b00001111110111100000000000000001;
mem[576] = 32'b00001111101000010000000000000000;
mem[577] = 32'b00110100000000010000000000111110;
mem[578] = 32'b00101100000000010000000000111110;
mem[579] = 32'b00101100000000100000000000111010;
mem[580] = 32'b00001000010000010000100000000000;
mem[581] = 32'b00101100001000010000000000000000;
mem[582] = 32'b00110100000000010000000000111111;
mem[583] = 32'b00101100000000010000000000111110;
mem[584] = 32'b00101100000000100000000000111010;
mem[585] = 32'b00001000010000010000100000000000;
mem[586] = 32'b00001100001001000000000000000000;
mem[587] = 32'b00101100000000010000000000111101;
mem[588] = 32'b00101100000000100000000000111010;
mem[589] = 32'b00001000010000010000100000000000;
mem[590] = 32'b00101100001000010000000000000000;
mem[591] = 32'b00110100100000010000000000000000;
mem[592] = 32'b00101100000000010000000000111101;
mem[593] = 32'b00101100000000100000000000111010;
mem[594] = 32'b00001000010000010000100000000000;
mem[595] = 32'b00001100001001000000000000000000;
mem[596] = 32'b00101100000000010000000000111111;
mem[597] = 32'b00110100100000010000000000000000;
mem[598] = 32'b00101100000000010000000000111101;
mem[599] = 32'b00001100001001000000000000000000;
mem[600] = 32'b00110000000000010000000000000001;
mem[601] = 32'b00001100001000100000000000000000;
mem[602] = 32'b00001100100000110000000000000000;
mem[603] = 32'b00001000011000100000100000000000;
mem[604] = 32'b00110100000000010000000000111101;
mem[605] = 32'b00111000000000000000001000100100;
mem[606] = 32'b00111111111000000000000000000000;
mem[607] = 32'b00110000000000010000000000000001;
mem[608] = 32'b00110100000000010000000001000000;
mem[609] = 32'b00101100000000010000000001000000;
mem[610] = 32'b00001100001001000000000000000000;
mem[611] = 32'b00110000000000010000000000000000;
mem[612] = 32'b00001100001000100000000000000000;
mem[613] = 32'b00001100100000110000000000000000;
mem[614] = 32'b01100000011000100000001011111011;
mem[615] = 32'b01111100000000010000000000000000;
mem[616] = 32'b00110100000000010000000001000000;
mem[617] = 32'b00101100000000010000000001000000;
mem[618] = 32'b00001100001001000000000000000000;
mem[619] = 32'b00110000000000010000000000000001;
mem[620] = 32'b00001100001000100000000000000000;
mem[621] = 32'b00001100100000110000000000000000;
mem[622] = 32'b01011100011000100000001001111100;
mem[623] = 32'b01111100000000010000000000000000;
mem[624] = 32'b00110100000000010000000001000011;
mem[625] = 32'b01111100000000010000000000000000;
mem[626] = 32'b00110100000000010000000001000100;
mem[627] = 32'b00101100000000010000000001000011;
mem[628] = 32'b00110100000000010000000000011011;
mem[629] = 32'b00101100000000010000000001000100;
mem[630] = 32'b00110100000000010000000000011100;
mem[631] = 32'b10000100000000000000000000110000;
mem[632] = 32'b00001111101000010000000000000000;
mem[633] = 32'b00110100000000010000000001000010;
mem[634] = 32'b10000000000000000000000001000010;
mem[635] = 32'b00111000000000000000001011111001;
mem[636] = 32'b00101100000000010000000001000000;
mem[637] = 32'b00001100001001000000000000000000;
mem[638] = 32'b00110000000000010000000000000010;
mem[639] = 32'b00001100001000100000000000000000;
mem[640] = 32'b00001100100000110000000000000000;
mem[641] = 32'b01011100011000100000001010001011;
mem[642] = 32'b01111100000000010000000000000000;
mem[643] = 32'b00110100000000010000000001000011;
mem[644] = 32'b00101100000000010000000001000011;
mem[645] = 32'b00110100000000010000000000110001;
mem[646] = 32'b10000100000000000000000110010001;
mem[647] = 32'b00001111101000010000000000000000;
mem[648] = 32'b00110100000000010000000001000010;
mem[649] = 32'b10000000000000000000000001000010;
mem[650] = 32'b00111000000000000000001011111001;
mem[651] = 32'b00101100000000010000000001000000;
mem[652] = 32'b00001100001001000000000000000000;
mem[653] = 32'b00110000000000010000000000000011;
mem[654] = 32'b00001100001000100000000000000000;
mem[655] = 32'b00001100100000110000000000000000;
mem[656] = 32'b01011100011000100000001010011010;
mem[657] = 32'b01111100000000010000000000000000;
mem[658] = 32'b00110100000000010000000001000011;
mem[659] = 32'b00101100000000010000000001000011;
mem[660] = 32'b00110100000000010000000000110000;
mem[661] = 32'b10000100000000000000000101011010;
mem[662] = 32'b00001111101000010000000000000000;
mem[663] = 32'b00110100000000010000000001000010;
mem[664] = 32'b10000000000000000000000001000010;
mem[665] = 32'b00111000000000000000001011111001;
mem[666] = 32'b00101100000000010000000001000000;
mem[667] = 32'b00001100001001000000000000000000;
mem[668] = 32'b00110000000000010000000000000100;
mem[669] = 32'b00001100001000100000000000000000;
mem[670] = 32'b00001100100000110000000000000000;
mem[671] = 32'b01011100011000100000001010110100;
mem[672] = 32'b01111100000000010000000000000000;
mem[673] = 32'b00110100000000010000000001000001;
mem[674] = 32'b00110000000000010000000000000000;
mem[675] = 32'b00110100000000010000000000010100;
mem[676] = 32'b00101100000000010000000001000001;
mem[677] = 32'b00110100000000010000000000010101;
mem[678] = 32'b10000100000000000000000000000010;
mem[679] = 32'b00110000000000010000000000000000;
mem[680] = 32'b00110100000000010000000000111010;
mem[681] = 32'b00110000000000010000000000000000;
mem[682] = 32'b00110100000000010000000000111011;
mem[683] = 32'b00101100000000010000000001000001;
mem[684] = 32'b00110100000000010000000000111100;
mem[685] = 32'b10000100000000000000001000100010;
mem[686] = 32'b00110000000000010000000000000000;
mem[687] = 32'b00110100000000010000000000010111;
mem[688] = 32'b00101100000000010000000001000001;
mem[689] = 32'b00110100000000010000000000011000;
mem[690] = 32'b10000100000000000000000000011001;
mem[691] = 32'b00111000000000000000001011111001;
mem[692] = 32'b00101100000000010000000001000000;
mem[693] = 32'b00001100001001000000000000000000;
mem[694] = 32'b00110000000000010000000000000101;
mem[695] = 32'b00001100001000100000000000000000;
mem[696] = 32'b00001100100000110000000000000000;
mem[697] = 32'b01011100011000100000001011000111;
mem[698] = 32'b01111100000000010000000000000000;
mem[699] = 32'b00110100000000010000000001000011;
mem[700] = 32'b01111100000000010000000000000000;
mem[701] = 32'b00110100000000010000000001000100;
mem[702] = 32'b00101100000000010000000001000011;
mem[703] = 32'b00110100000000010000000000110010;
mem[704] = 32'b00101100000000010000000001000100;
mem[705] = 32'b00110100000000010000000000110011;
mem[706] = 32'b10000100000000000000000111000000;
mem[707] = 32'b00001111101000010000000000000000;
mem[708] = 32'b00110100000000010000000001000010;
mem[709] = 32'b10000000000000000000000001000010;
mem[710] = 32'b00111000000000000000001011111001;
mem[711] = 32'b00101100000000010000000001000000;
mem[712] = 32'b00001100001001000000000000000000;
mem[713] = 32'b00110000000000010000000000000110;
mem[714] = 32'b00001100001000100000000000000000;
mem[715] = 32'b00001100100000110000000000000000;
mem[716] = 32'b01011100011000100000001011100101;
mem[717] = 32'b01111100000000010000000000000000;
mem[718] = 32'b00110100000000010000000001000001;
mem[719] = 32'b00110000000000010000000000000000;
mem[720] = 32'b00110100000000010000000000010100;
mem[721] = 32'b00101100000000010000000001000001;
mem[722] = 32'b00110100000000010000000000010101;
mem[723] = 32'b10000100000000000000000000000010;
mem[724] = 32'b00110000000000010000000000000000;
mem[725] = 32'b00110100000000010000000000101100;
mem[726] = 32'b00101100000000010000000001000001;
mem[727] = 32'b00110100000000010000000000101101;
mem[728] = 32'b10000100000000000000000100110100;
mem[729] = 32'b00001111101000010000000000000000;
mem[730] = 32'b00110100000000010000000001000010;
mem[731] = 32'b10000000000000000000000001000010;
mem[732] = 32'b00110000000000010000000000000000;
mem[733] = 32'b00110100000000010000000000101000;
mem[734] = 32'b00101100000000010000000001000001;
mem[735] = 32'b00110100000000010000000000101001;
mem[736] = 32'b10000100000000000000000100001110;
mem[737] = 32'b00001111101000010000000000000000;
mem[738] = 32'b00110100000000010000000001000010;
mem[739] = 32'b10000000000000000000000001000010;
mem[740] = 32'b00111000000000000000001011111001;
mem[741] = 32'b00101100000000010000000001000000;
mem[742] = 32'b00001100001001000000000000000000;
mem[743] = 32'b00110000000000010000000000000111;
mem[744] = 32'b00001100001000100000000000000000;
mem[745] = 32'b00001100100000110000000000000000;
mem[746] = 32'b01011100011000100000001011111010;
mem[747] = 32'b01111100000000010000000000000000;
mem[748] = 32'b00110100000000010000000001000001;
mem[749] = 32'b00110000000000010000000000000000;
mem[750] = 32'b00110100000000010000000000010100;
mem[751] = 32'b00101100000000010000000001000001;
mem[752] = 32'b00110100000000010000000000010101;
mem[753] = 32'b10000100000000000000000000000010;
mem[754] = 32'b00110000000000010000000000000000;
mem[755] = 32'b00110100000000010000000000011111;
mem[756] = 32'b00101100000000010000000001000001;
mem[757] = 32'b00110100000000010000000000100000;
mem[758] = 32'b10000100000000000000000001001100;
mem[759] = 32'b00001111101000010000000000000000;
mem[760] = 32'b00110100000000010000000001000010;
mem[761] = 32'b10000000000000000000000001000010;
mem[762] = 32'b00111000000000000000001001100001;
mem[763] = 32'b00000100000000000000000000000000;
			end
		end
	always @( posedge autoclock )
		begin
			InstructionOut = mem[adress];
		end
endmodule
	
