module InstructionMemory #(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=1900, parameter TRACKS=2)
(address, InstructionOut, clock, autoclock, rst, writeInstr, instrIn, pId, WritepId, HDAddress, region );

	input [(DATA_WIDTH-1):0] address, HDAddress, pId, WritepId, instrIn;
	input clock, autoclock, rst, writeInstr;
	input region;
	output reg [(DATA_WIDTH-1):0] InstructionOut;
	reg [(DATA_WIDTH-1):0] mem [((ADDR_WIDTH*TRACKS)-1):0];
	
	initial begin
/*mem[0] = 32'b00000000000000000000000000000000;
mem[1] = 32'b00111000000000000000010100011100;
mem[2] = 32'b00110000000000010000000000000000;
mem[3] = 32'b00001100001001000000000000000000;
mem[4] = 32'b00110000000000010000000000000000;
mem[5] = 32'b00110100100000010000000000000100;
mem[6] = 32'b00110000000000010000000000000000;
mem[7] = 32'b00001100001001000000000000000000;
mem[8] = 32'b00110000000000010000000000000000;
mem[9] = 32'b00110100100000010000000000100111;
mem[10] = 32'b00110000000000010000000000000000;
mem[11] = 32'b00001100001001000000000000000000;
mem[12] = 32'b00110000000000010000011101010111;
mem[13] = 32'b00110100100000010000000001001010;
mem[14] = 32'b00110000000000010000000000000000;
mem[15] = 32'b00001100001001000000000000000000;
mem[16] = 32'b00110000000000010000000000000000;
mem[17] = 32'b00110100100000010000000001101101;
mem[18] = 32'b00110000000000010000000000000000;
mem[19] = 32'b00001100001001000000000000000000;
mem[20] = 32'b00110000000000010000000000000001;
mem[21] = 32'b00110100100000010000000010010000;
mem[22] = 32'b00110000000000010000000000000000;
mem[23] = 32'b00001100001001000000000000000000;
mem[24] = 32'b00110000000000010000011101011000;
mem[25] = 32'b00110100100000010000000010110011;
mem[26] = 32'b00110000000000010000000000000001;
mem[27] = 32'b00110100000000010000000011010110;
mem[28] = 32'b00110000000000010000000000000001;
mem[29] = 32'b00110100000000010000000011010111;
mem[30] = 32'b00110000000000010000000000000001;
mem[31] = 32'b00110100000000010000000100001010;
mem[32] = 32'b00110000000000010000011101011000;
mem[33] = 32'b00110100000000010000000100001011;
mem[34] = 32'b00110000000000010000000000100000;
mem[35] = 32'b00110100000000010000000100001100;
mem[36] = 32'b00101100000000010000000011010110;
mem[37] = 32'b00110100000000010000000011011000;
mem[38] = 32'b00101100000000010000000011010110;
mem[39] = 32'b00001100001001000000000000000000;
mem[40] = 32'b00110000000000010000000000000001;
mem[41] = 32'b00110100100000010000000000000100;
mem[42] = 32'b00101100000000010000000011010110;
mem[43] = 32'b00001100001001000000000000000000;
mem[44] = 32'b00110000000000010000000000000000;
mem[45] = 32'b00110100100000010000000000100111;
mem[46] = 32'b00101100000000010000000011010110;
mem[47] = 32'b00001100001001000000000000000000;
mem[48] = 32'b00110000000000010000000000001000;
mem[49] = 32'b00110100100000010000000001001010;
mem[50] = 32'b00101100000000010000000011010110;
mem[51] = 32'b00001100001001000000000000000000;
mem[52] = 32'b00110000000000010000000000110010;
mem[53] = 32'b00110100100000010000000001101101;
mem[54] = 32'b00101100000000010000000011010110;
mem[55] = 32'b00001100001001000000000000000000;
mem[56] = 32'b00110000000000010000000000000001;
mem[57] = 32'b00110100100000010000000010010000;
mem[58] = 32'b00101100000000010000000011010110;
mem[59] = 32'b00001100001001000000000000000000;
mem[60] = 32'b00110000000000010000000000001001;
mem[61] = 32'b00110100100000010000000010110011;
mem[62] = 32'b00101100000000010000000011010110;
mem[63] = 32'b00001100001001000000000000000000;
mem[64] = 32'b00110000000000010000000000000001;
mem[65] = 32'b00001100001000100000000000000000;
mem[66] = 32'b00001100100000110000000000000000;
mem[67] = 32'b00001000011000100000100000000000;
mem[68] = 32'b00110100000000010000000011010110;
mem[69] = 32'b00101100000000010000000011010110;
mem[70] = 32'b00001100001001000000000000000000;
mem[71] = 32'b00110000000000010000000000000001;
mem[72] = 32'b00110100100000010000000000000100;
mem[73] = 32'b00101100000000010000000011010110;
mem[74] = 32'b00001100001001000000000000000000;
mem[75] = 32'b00110000000000010000000001001101;
mem[76] = 32'b00110100100000010000000000100111;
mem[77] = 32'b00101100000000010000000011010110;
mem[78] = 32'b00001100001001000000000000000000;
mem[79] = 32'b00110000000000010000000010001111;
mem[80] = 32'b00110100100000010000000001001010;
mem[81] = 32'b00101100000000010000000011010110;
mem[82] = 32'b00001100001001000000000000000000;
mem[83] = 32'b00110000000000010000000000110011;
mem[84] = 32'b00110100100000010000000001101101;
mem[85] = 32'b00101100000000010000000011010110;
mem[86] = 32'b00001100001001000000000000000000;
mem[87] = 32'b00110000000000010000000000000001;
mem[88] = 32'b00110100100000010000000010010000;
mem[89] = 32'b00101100000000010000000011010110;
mem[90] = 32'b00001100001001000000000000000000;
mem[91] = 32'b00110000000000010000000001000011;
mem[92] = 32'b00110100100000010000000010110011;
mem[93] = 32'b00101100000000010000000011010110;
mem[94] = 32'b00001100001001000000000000000000;
mem[95] = 32'b00110000000000010000000000000001;
mem[96] = 32'b00001100001000100000000000000000;
mem[97] = 32'b00001100100000110000000000000000;
mem[98] = 32'b00001000011000100000100000000000;
mem[99] = 32'b00110100000000010000000011010110;
mem[100] = 32'b00101100000000010000000011010110;
mem[101] = 32'b00001100001001000000000000000000;
mem[102] = 32'b00110000000000010000000000000001;
mem[103] = 32'b00110100100000010000000000000100;
mem[104] = 32'b00101100000000010000000011010110;
mem[105] = 32'b00001100001001000000000000000000;
mem[106] = 32'b00110000000000010000000010010000;
mem[107] = 32'b00110100100000010000000000100111;
mem[108] = 32'b00101100000000010000000011010110;
mem[109] = 32'b00001100001001000000000000000000;
mem[110] = 32'b00110000000000010000000011000011;
mem[111] = 32'b00110100100000010000000001001010;
mem[112] = 32'b00101100000000010000000011010110;
mem[113] = 32'b00001100001001000000000000000000;
mem[114] = 32'b00110000000000010000000000110100;
mem[115] = 32'b00110100100000010000000001101101;
mem[116] = 32'b00101100000000010000000011010110;
mem[117] = 32'b00001100001001000000000000000000;
mem[118] = 32'b00110000000000010000000000000001;
mem[119] = 32'b00110100100000010000000010010000;
mem[120] = 32'b00101100000000010000000011010110;
mem[121] = 32'b00001100001001000000000000000000;
mem[122] = 32'b00110000000000010000000000110100;
mem[123] = 32'b00110100100000010000000010110011;
mem[124] = 32'b00101100000000010000000011010110;
mem[125] = 32'b00001100001001000000000000000000;
mem[126] = 32'b00110000000000010000000000000001;
mem[127] = 32'b00001100001000100000000000000000;
mem[128] = 32'b00001100100000110000000000000000;
mem[129] = 32'b00001000011000100000100000000000;
mem[130] = 32'b00110100000000010000000011010110;
mem[131] = 32'b00101100000000010000000011010110;
mem[132] = 32'b00001100001001000000000000000000;
mem[133] = 32'b00110000000000010000000000000001;
mem[134] = 32'b00110100100000010000000000000100;
mem[135] = 32'b00101100000000010000000011010110;
mem[136] = 32'b00001100001001000000000000000000;
mem[137] = 32'b00110000000000010000000011000100;
mem[138] = 32'b00110100100000010000000000100111;
mem[139] = 32'b00101100000000010000000011010110;
mem[140] = 32'b00001100001001000000000000000000;
mem[141] = 32'b00110000000000010000000100011111;
mem[142] = 32'b00110100100000010000000001001010;
mem[143] = 32'b00101100000000010000000011010110;
mem[144] = 32'b00001100001001000000000000000000;
mem[145] = 32'b00110000000000010000000000110101;
mem[146] = 32'b00110100100000010000000001101101;
mem[147] = 32'b00101100000000010000000011010110;
mem[148] = 32'b00001100001001000000000000000000;
mem[149] = 32'b00110000000000010000000000000001;
mem[150] = 32'b00110100100000010000000010010000;
mem[151] = 32'b00101100000000010000000011010110;
mem[152] = 32'b00001100001001000000000000000000;
mem[153] = 32'b00110000000000010000000001011100;
mem[154] = 32'b00110100100000010000000010110011;
mem[155] = 32'b00101100000000010000000011010110;
mem[156] = 32'b00001100001001000000000000000000;
mem[157] = 32'b00110000000000010000000000000001;
mem[158] = 32'b00001100001000100000000000000000;
mem[159] = 32'b00001100100000110000000000000000;
mem[160] = 32'b00001000011000100000100000000000;
mem[161] = 32'b00110100000000010000000011010110;
mem[162] = 32'b00101100000000010000000011010110;
mem[163] = 32'b00001100001001000000000000000000;
mem[164] = 32'b00110000000000010000000000000001;
mem[165] = 32'b00110100100000010000000000000100;
mem[166] = 32'b00101100000000010000000011010110;
mem[167] = 32'b00001100001001000000000000000000;
mem[168] = 32'b00110000000000010000000100100000;
mem[169] = 32'b00110100100000010000000000100111;
mem[170] = 32'b00101100000000010000000011010110;
mem[171] = 32'b00001100001001000000000000000000;
mem[172] = 32'b00110000000000010000000101111101;
mem[173] = 32'b00110100100000010000000001001010;
mem[174] = 32'b00101100000000010000000011010110;
mem[175] = 32'b00001100001001000000000000000000;
mem[176] = 32'b00110000000000010000000000110110;
mem[177] = 32'b00110100100000010000000001101101;
mem[178] = 32'b00101100000000010000000011010110;
mem[179] = 32'b00001100001001000000000000000000;
mem[180] = 32'b00110000000000010000000000000001;
mem[181] = 32'b00110100100000010000000010010000;
mem[182] = 32'b00101100000000010000000011010110;
mem[183] = 32'b00001100001001000000000000000000;
mem[184] = 32'b00110000000000010000000001011110;
mem[185] = 32'b00110100100000010000000010110011;
mem[186] = 32'b00101100000000010000000011010110;
mem[187] = 32'b00001100001001000000000000000000;
mem[188] = 32'b00110000000000010000000000000001;
mem[189] = 32'b00001100001000100000000000000000;
mem[190] = 32'b00001100100000110000000000000000;
mem[191] = 32'b00001000011000100000100000000000;
mem[192] = 32'b00110100000000010000000011010110;
mem[193] = 32'b00101100000000010000000011010110;
mem[194] = 32'b00001100001001000000000000000000;
mem[195] = 32'b00110000000000010000000000000001;
mem[196] = 32'b00110100100000010000000000000100;
mem[197] = 32'b00101100000000010000000011010110;
mem[198] = 32'b00001100001001000000000000000000;
mem[199] = 32'b00110000000000010000000101111110;
mem[200] = 32'b00110100100000010000000000100111;
mem[201] = 32'b00101100000000010000000011010110;
mem[202] = 32'b00001100001001000000000000000000;
mem[203] = 32'b00110000000000010000000111011011;
mem[204] = 32'b00110100100000010000000001001010;
mem[205] = 32'b00101100000000010000000011010110;
mem[206] = 32'b00001100001001000000000000000000;
mem[207] = 32'b00110000000000010000000000110111;
mem[208] = 32'b00110100100000010000000001101101;
mem[209] = 32'b00101100000000010000000011010110;
mem[210] = 32'b00001100001001000000000000000000;
mem[211] = 32'b00110000000000010000000000000001;
mem[212] = 32'b00110100100000010000000010010000;
mem[213] = 32'b00101100000000010000000011010110;
mem[214] = 32'b00001100001001000000000000000000;
mem[215] = 32'b00110000000000010000000001011110;
mem[216] = 32'b00110100100000010000000010110011;
mem[217] = 32'b00101100000000010000000011010110;
mem[218] = 32'b00001100001001000000000000000000;
mem[219] = 32'b00110000000000010000000000000001;
mem[220] = 32'b00001100001000100000000000000000;
mem[221] = 32'b00001100100000110000000000000000;
mem[222] = 32'b00001000011000100000100000000000;
mem[223] = 32'b00110100000000010000000011010110;
mem[224] = 32'b00101100000000010000000011010110;
mem[225] = 32'b00001100001001000000000000000000;
mem[226] = 32'b00110000000000010000000000000001;
mem[227] = 32'b00110100100000010000000000000100;
mem[228] = 32'b00101100000000010000000011010110;
mem[229] = 32'b00001100001001000000000000000000;
mem[230] = 32'b00110000000000010000000111011100;
mem[231] = 32'b00110100100000010000000000100111;
mem[232] = 32'b00101100000000010000000011010110;
mem[233] = 32'b00001100001001000000000000000000;
mem[234] = 32'b00110000000000010000001000101000;
mem[235] = 32'b00110100100000010000000001001010;
mem[236] = 32'b00101100000000010000000011010110;
mem[237] = 32'b00001100001001000000000000000000;
mem[238] = 32'b00110000000000010000000000111000;
mem[239] = 32'b00110100100000010000000001101101;
mem[240] = 32'b00101100000000010000000011010110;
mem[241] = 32'b00001100001001000000000000000000;
mem[242] = 32'b00110000000000010000000000000001;
mem[243] = 32'b00110100100000010000000010010000;
mem[244] = 32'b00101100000000010000000011010110;
mem[245] = 32'b00001100001001000000000000000000;
mem[246] = 32'b00110000000000010000000001001101;
mem[247] = 32'b00110100100000010000000010110011;
mem[248] = 32'b00101100000000010000000011010110;
mem[249] = 32'b00001100001001000000000000000000;
mem[250] = 32'b00110000000000010000000000000001;
mem[251] = 32'b00001100001000100000000000000000;
mem[252] = 32'b00001100100000110000000000000000;
mem[253] = 32'b00001000011000100000100000000000;
mem[254] = 32'b00110100000000010000000011010110;
mem[255] = 32'b00101100000000010000000011010110;
mem[256] = 32'b00001100001001000000000000000000;
mem[257] = 32'b00110000000000010000000000000001;
mem[258] = 32'b00110100100000010000000000000100;
mem[259] = 32'b00101100000000010000000011010110;
mem[260] = 32'b00001100001001000000000000000000;
mem[261] = 32'b00110000000000010000001000101001;
mem[262] = 32'b00110100100000010000000000100111;
mem[263] = 32'b00101100000000010000000011010110;
mem[264] = 32'b00001100001001000000000000000000;
mem[265] = 32'b00110000000000010000001001110011;
mem[266] = 32'b00110100100000010000000001001010;
mem[267] = 32'b00101100000000010000000011010110;
mem[268] = 32'b00001100001001000000000000000000;
mem[269] = 32'b00110000000000010000000000111001;
mem[270] = 32'b00110100100000010000000001101101;
mem[271] = 32'b00101100000000010000000011010110;
mem[272] = 32'b00001100001001000000000000000000;
mem[273] = 32'b00110000000000010000000000000001;
mem[274] = 32'b00110100100000010000000010010000;
mem[275] = 32'b00101100000000010000000011010110;
mem[276] = 32'b00001100001001000000000000000000;
mem[277] = 32'b00110000000000010000000001001011;
mem[278] = 32'b00110100100000010000000010110011;
mem[279] = 32'b00101100000000010000000011010110;
mem[280] = 32'b00001100001001000000000000000000;
mem[281] = 32'b00110000000000010000000000000001;
mem[282] = 32'b00001100001000100000000000000000;
mem[283] = 32'b00001100100000110000000000000000;
mem[284] = 32'b00001000011000100000100000000000;
mem[285] = 32'b00110100000000010000000011010110;
mem[286] = 32'b00101100000000010000000011010110;
mem[287] = 32'b00001100001001000000000000000000;
mem[288] = 32'b00110000000000010000000000000001;
mem[289] = 32'b00110100100000010000000000000100;
mem[290] = 32'b00101100000000010000000011010110;
mem[291] = 32'b00001100001001000000000000000000;
mem[292] = 32'b00110000000000010000001001110100;
mem[293] = 32'b00110100100000010000000000100111;
mem[294] = 32'b00101100000000010000000011010110;
mem[295] = 32'b00001100001001000000000000000000;
mem[296] = 32'b00110000000000010000001011010010;
mem[297] = 32'b00110100100000010000000001001010;
mem[298] = 32'b00101100000000010000000011010110;
mem[299] = 32'b00001100001001000000000000000000;
mem[300] = 32'b00110000000000010000000000111010;
mem[301] = 32'b00110100100000010000000001101101;
mem[302] = 32'b00101100000000010000000011010110;
mem[303] = 32'b00001100001001000000000000000000;
mem[304] = 32'b00110000000000010000000000000001;
mem[305] = 32'b00110100100000010000000010010000;
mem[306] = 32'b00101100000000010000000011010110;
mem[307] = 32'b00001100001001000000000000000000;
mem[308] = 32'b00110000000000010000000001011111;
mem[309] = 32'b00110100100000010000000010110011;
mem[310] = 32'b00101100000000010000000011010110;
mem[311] = 32'b00001100001001000000000000000000;
mem[312] = 32'b00110000000000010000000000000001;
mem[313] = 32'b00001100001000100000000000000000;
mem[314] = 32'b00001100100000110000000000000000;
mem[315] = 32'b00001000011000100000100000000000;
mem[316] = 32'b00110100000000010000000011010110;
mem[317] = 32'b00101100000000010000000011010110;
mem[318] = 32'b00001100001001000000000000000000;
mem[319] = 32'b00110000000000010000000000000001;
mem[320] = 32'b00110100100000010000000000000100;
mem[321] = 32'b00101100000000010000000011010110;
mem[322] = 32'b00001100001001000000000000000000;
mem[323] = 32'b00110000000000010000001011010011;
mem[324] = 32'b00110100100000010000000000100111;
mem[325] = 32'b00101100000000010000000011010110;
mem[326] = 32'b00001100001001000000000000000000;
mem[327] = 32'b00110000000000010000001100000010;
mem[328] = 32'b00110100100000010000000001001010;
mem[329] = 32'b00101100000000010000000011010110;
mem[330] = 32'b00001100001001000000000000000000;
mem[331] = 32'b00110000000000010000000000111011;
mem[332] = 32'b00110100100000010000000001101101;
mem[333] = 32'b00101100000000010000000011010110;
mem[334] = 32'b00001100001001000000000000000000;
mem[335] = 32'b00110000000000010000000000000001;
mem[336] = 32'b00110100100000010000000010010000;
mem[337] = 32'b00101100000000010000000011010110;
mem[338] = 32'b00001100001001000000000000000000;
mem[339] = 32'b00110000000000010000000000110000;
mem[340] = 32'b00110100100000010000000010110011;
mem[341] = 32'b00101100000000010000000011010110;
mem[342] = 32'b00001100001001000000000000000000;
mem[343] = 32'b00110000000000010000000000000001;
mem[344] = 32'b00001100001000100000000000000000;
mem[345] = 32'b00001100100000110000000000000000;
mem[346] = 32'b00001000011000100000100000000000;
mem[347] = 32'b00110100000000010000000011010110;
mem[348] = 32'b00111111111000000000000000000000;
mem[349] = 32'b00110000000000010000000000000001;
mem[350] = 32'b00110100000000010000000011111011;
mem[351] = 32'b00110000000000010000000000000010;
mem[352] = 32'b00110100000000010000000011111100;
mem[353] = 32'b00110000000000010000000000000011;
mem[354] = 32'b00110100000000010000000011111101;
mem[355] = 32'b00110000000000010000000000000100;
mem[356] = 32'b00110100000000010000000011111110;
mem[357] = 32'b00110000000000010000000000000101;
mem[358] = 32'b00110100000000010000000011111111;
mem[359] = 32'b00110000000000010000000000000110;
mem[360] = 32'b00110100000000010000000100000000;
mem[361] = 32'b00110000000000010000000000000111;
mem[362] = 32'b00110100000000010000000100000001;
mem[363] = 32'b00110000000000010000000000001000;
mem[364] = 32'b00110100000000010000000100000010;
mem[365] = 32'b00110000000000010000000000001001;
mem[366] = 32'b00110100000000010000000100000011;
mem[367] = 32'b00110000000000010000000000001010;
mem[368] = 32'b00110100000000010000000100000100;
mem[369] = 32'b00110000000000010000000000001011;
mem[370] = 32'b00110100000000010000000100000101;
mem[371] = 32'b00110000000000010000000000001100;
mem[372] = 32'b00110100000000010000000100000110;
mem[373] = 32'b00110000000000010000011111001111;
mem[374] = 32'b00110100000000010000000100000111;
mem[375] = 32'b00110000000000010000000000000101;
mem[376] = 32'b00110100000000010000000100001000;
mem[377] = 32'b00101100000000010000000011111011;
mem[378] = 32'b10011000001000000000000000000000;
mem[379] = 32'b00001111110111101111111111111111;
mem[380] = 32'b00110111110111110000000000000000;
mem[381] = 32'b10000100000000000000000000000010;
mem[382] = 32'b00101111110111110000000000000000;
mem[383] = 32'b00001111110111100000000000000001;
mem[384] = 32'b00111111111000000000000000000000;
mem[385] = 32'b00111111111000000000000000000000;
mem[386] = 32'b00110000000000010000000000000000;
mem[387] = 32'b00110100000000010000000100001110;
mem[388] = 32'b00101100000000010000000100001110;
mem[389] = 32'b00001100001001000000000000000000;
mem[390] = 32'b00101100000000010000000011010110;
mem[391] = 32'b00001100001000100000000000000000;
mem[392] = 32'b00001100100000110000000000000000;
mem[393] = 32'b01110000011000100000000110011100;
mem[394] = 32'b00101100000000010000000100001110;
mem[395] = 32'b00101100001000010000000001101101;
mem[396] = 32'b00001100001001000000000000000000;
mem[397] = 32'b00101100000000010000000100001101;
mem[398] = 32'b00001100001000100000000000000000;
mem[399] = 32'b00001100100000110000000000000000;
mem[400] = 32'b01011100011000100000000110010100;
mem[401] = 32'b00101100000000010000000100001110;
mem[402] = 32'b00001100001111010000000000000000;
mem[403] = 32'b00111111111000000000000000000000;
mem[404] = 32'b00101100000000010000000100001110;
mem[405] = 32'b00001100001001000000000000000000;
mem[406] = 32'b00110000000000010000000000000001;
mem[407] = 32'b00001100001000100000000000000000;
mem[408] = 32'b00001100100000110000000000000000;
mem[409] = 32'b00001000011000100000100000000000;
mem[410] = 32'b00110100000000010000000100001110;
mem[411] = 32'b00111000000000000000000110000100;
mem[412] = 32'b00110000000000010000000000000000;
mem[413] = 32'b00001100001111010000000000000000;
mem[414] = 32'b00111111111000000000000000000000;
mem[415] = 32'b00110000000000010000000000000000;
mem[416] = 32'b00110100000000010000000100010000;
mem[417] = 32'b00110000000000010000000001100011;
mem[418] = 32'b00110100000000010000000100010001;
mem[419] = 32'b00101100000000010000000011111111;
mem[420] = 32'b10011000001000000000000000000000;
mem[421] = 32'b01111100000000010000000000000000;
mem[422] = 32'b00110100000000010000000100010010;
mem[423] = 32'b01111100000000010000000000000000;
mem[424] = 32'b00110100000000010000000100010011;
mem[425] = 32'b00101100000000010000000100010000;
mem[426] = 32'b00001100001001000000000000000000;
mem[427] = 32'b00101100000000010000000011010110;
mem[428] = 32'b00001100001000100000000000000000;
mem[429] = 32'b00001100100000110000000000000000;
mem[430] = 32'b01110000011000100000000111001100;
mem[431] = 32'b00101100000000010000000100010000;
mem[432] = 32'b00101100001000010000000010010000;
mem[433] = 32'b00001100001001000000000000000000;
mem[434] = 32'b00110000000000010000000000000000;
mem[435] = 32'b00001100001000100000000000000000;
mem[436] = 32'b00001100100000110000000000000000;
mem[437] = 32'b01011100011000100000000110111001;
mem[438] = 32'b00110000000000010000000001100011;
mem[439] = 32'b00110100000000010000000100010000;
mem[440] = 32'b00111000000000000000000111000100;
mem[441] = 32'b00101100000000010000000100010000;
mem[442] = 32'b00101100001000010000000001101101;
mem[443] = 32'b00001100001001000000000000000000;
mem[444] = 32'b00101100000000010000000100010010;
mem[445] = 32'b00001100001000100000000000000000;
mem[446] = 32'b00001100100000110000000000000000;
mem[447] = 32'b01011100011000100000000111000100;
mem[448] = 32'b00101100000000010000000100010000;
mem[449] = 32'b00110100000000010000000100010001;
mem[450] = 32'b00110000000000010000000001100011;
mem[451] = 32'b00110100000000010000000100010000;
mem[452] = 32'b00101100000000010000000100010000;
mem[453] = 32'b00001100001001000000000000000000;
mem[454] = 32'b00110000000000010000000000000001;
mem[455] = 32'b00001100001000100000000000000000;
mem[456] = 32'b00001100100000110000000000000000;
mem[457] = 32'b00001000011000100000100000000000;
mem[458] = 32'b00110100000000010000000100010000;
mem[459] = 32'b00111000000000000000000110101001;
mem[460] = 32'b00101100000000010000000100010001;
mem[461] = 32'b00001100001001000000000000000000;
mem[462] = 32'b00101100000000010000000011010110;
mem[463] = 32'b00001100001000100000000000000000;
mem[464] = 32'b00001100100000110000000000000000;
mem[465] = 32'b01110000011000100000000111010110;
mem[466] = 32'b00101100000000010000000100010001;
mem[467] = 32'b00001100001001000000000000000000;
mem[468] = 32'b00101100000000010000000100010011;
mem[469] = 32'b00110100100000010000000001101101;
mem[470] = 32'b00111111111000000000000000000000;
mem[471] = 32'b00101100000000010000000100000000;
mem[472] = 32'b10011000001000000000000000000000;
mem[473] = 32'b01111100000000010000000000000000;
mem[474] = 32'b00110100000000010000000000000011;
mem[475] = 32'b00101100000000010000000011011000;
mem[476] = 32'b00110100000000010000000100010100;
mem[477] = 32'b00110000000000010000000000000001;
mem[478] = 32'b00110100000000010000000100010101;
mem[479] = 32'b00101100000000010000000100010101;
mem[480] = 32'b00001100001001000000000000000000;
mem[481] = 32'b00110000000000010000000000000000;
mem[482] = 32'b00001100001000100000000000000000;
mem[483] = 32'b00001100100000110000000000000000;
mem[484] = 32'b01100000011000100000001001100001;
mem[485] = 32'b00101100000000010000000100010100;
mem[486] = 32'b00101100001000010000000010010000;
mem[487] = 32'b00001100001001000000000000000000;
mem[488] = 32'b00110000000000010000000000000000;
mem[489] = 32'b00001100001000100000000000000000;
mem[490] = 32'b00001100100000110000000000000000;
mem[491] = 32'b01011100011000100000000111101111;
mem[492] = 32'b00110000000000010000000000000000;
mem[493] = 32'b00110100000000010000000100010101;
mem[494] = 32'b00111000000000000000001001100000;
mem[495] = 32'b00101100000000010000000100010100;
mem[496] = 32'b00101100001000010000000001101101;
mem[497] = 32'b00001100001001000000000000000000;
mem[498] = 32'b00101100000000010000000000000011;
mem[499] = 32'b00001100001000100000000000000000;
mem[500] = 32'b00001100100000110000000000000000;
mem[501] = 32'b01011100011000100000001001011001;
mem[502] = 32'b00101100000000010000000100010100;
mem[503] = 32'b00001100001001000000000000000000;
mem[504] = 32'b00110000000000010000000000000000;
mem[505] = 32'b00110100100000010000000010010000;
mem[506] = 32'b00110000000000010000000000000000;
mem[507] = 32'b00110100000000010000000100010101;
mem[508] = 32'b00101100000000010000000011010110;
mem[509] = 32'b00001100001001000000000000000000;
mem[510] = 32'b00101100000000010000000100010100;
mem[511] = 32'b00001100001000100000000000000000;
mem[512] = 32'b00001100100000110000000000000000;
mem[513] = 32'b01100000011000100000001001011001;
mem[514] = 32'b00101100000000010000000100010100;
mem[515] = 32'b00001100001001000000000000000000;
mem[516] = 32'b00110000000000010000000000000001;
mem[517] = 32'b00001100001000100000000000000000;
mem[518] = 32'b00001100100000110000000000000000;
mem[519] = 32'b00001000011000100000100000000000;
mem[520] = 32'b00101100001000010000000010010000;
mem[521] = 32'b00001100001001000000000000000000;
mem[522] = 32'b00110000000000010000000000000000;
mem[523] = 32'b00001100001000100000000000000000;
mem[524] = 32'b00001100100000110000000000000000;
mem[525] = 32'b01100000011000100000001001010010;
mem[526] = 32'b00101100000000010000000100010100;
mem[527] = 32'b00001100001001000000000000000000;
mem[528] = 32'b00101100000000010000000100010100;
mem[529] = 32'b00001100001001010000000000000000;
mem[530] = 32'b00110000000000010000000000000001;
mem[531] = 32'b00001100001000100000000000000000;
mem[532] = 32'b00001100101000110000000000000000;
mem[533] = 32'b00001000011000100000100000000000;
mem[534] = 32'b00101100001000010000000000000100;
mem[535] = 32'b00110100100000010000000000000100;
mem[536] = 32'b00101100000000010000000100010100;
mem[537] = 32'b00001100001001000000000000000000;
mem[538] = 32'b00101100000000010000000100010100;
mem[539] = 32'b00001100001001010000000000000000;
mem[540] = 32'b00110000000000010000000000000001;
mem[541] = 32'b00001100001000100000000000000000;
mem[542] = 32'b00001100101000110000000000000000;
mem[543] = 32'b00001000011000100000100000000000;
mem[544] = 32'b00101100001000010000000000100111;
mem[545] = 32'b00110100100000010000000000100111;
mem[546] = 32'b00101100000000010000000100010100;
mem[547] = 32'b00001100001001000000000000000000;
mem[548] = 32'b00101100000000010000000100010100;
mem[549] = 32'b00001100001001010000000000000000;
mem[550] = 32'b00110000000000010000000000000001;
mem[551] = 32'b00001100001000100000000000000000;
mem[552] = 32'b00001100101000110000000000000000;
mem[553] = 32'b00001000011000100000100000000000;
mem[554] = 32'b00101100001000010000000001001010;
mem[555] = 32'b00110100100000010000000001001010;
mem[556] = 32'b00101100000000010000000100010100;
mem[557] = 32'b00001100001001000000000000000000;
mem[558] = 32'b00101100000000010000000100010100;
mem[559] = 32'b00001100001001010000000000000000;
mem[560] = 32'b00110000000000010000000000000001;
mem[561] = 32'b00001100001000100000000000000000;
mem[562] = 32'b00001100101000110000000000000000;
mem[563] = 32'b00001000011000100000100000000000;
mem[564] = 32'b00101100001000010000000001101101;
mem[565] = 32'b00110100100000010000000001101101;
mem[566] = 32'b00101100000000010000000100010100;
mem[567] = 32'b00001100001001000000000000000000;
mem[568] = 32'b00101100000000010000000100010100;
mem[569] = 32'b00001100001001010000000000000000;
mem[570] = 32'b00110000000000010000000000000001;
mem[571] = 32'b00001100001000100000000000000000;
mem[572] = 32'b00001100101000110000000000000000;
mem[573] = 32'b00001000011000100000100000000000;
mem[574] = 32'b00101100001000010000000010010000;
mem[575] = 32'b00110100100000010000000010010000;
mem[576] = 32'b00101100000000010000000100010100;
mem[577] = 32'b00001100001001000000000000000000;
mem[578] = 32'b00101100000000010000000100010100;
mem[579] = 32'b00001100001001010000000000000000;
mem[580] = 32'b00110000000000010000000000000001;
mem[581] = 32'b00001100001000100000000000000000;
mem[582] = 32'b00001100101000110000000000000000;
mem[583] = 32'b00001000011000100000100000000000;
mem[584] = 32'b00101100001000010000000010110011;
mem[585] = 32'b00110100100000010000000010110011;
mem[586] = 32'b00101100000000010000000100010100;
mem[587] = 32'b00001100001001000000000000000000;
mem[588] = 32'b00110000000000010000000000000001;
mem[589] = 32'b00001100001000100000000000000000;
mem[590] = 32'b00001100100000110000000000000000;
mem[591] = 32'b00001000011000100000100000000000;
mem[592] = 32'b00110100000000010000000100010100;
mem[593] = 32'b00111000000000000000001000000010;
mem[594] = 32'b00101100000000010000000011010110;
mem[595] = 32'b00001100001001000000000000000000;
mem[596] = 32'b00110000000000010000000000000001;
mem[597] = 32'b00001100001000100000000000000000;
mem[598] = 32'b00001100100000110000000000000000;
mem[599] = 32'b00010000011000100000100000000000;
mem[600] = 32'b00110100000000010000000011010110;
mem[601] = 32'b00101100000000010000000100010100;
mem[602] = 32'b00001100001001000000000000000000;
mem[603] = 32'b00110000000000010000000000000001;
mem[604] = 32'b00001100001000100000000000000000;
mem[605] = 32'b00001100100000110000000000000000;
mem[606] = 32'b00001000011000100000100000000000;
mem[607] = 32'b00110100000000010000000100010100;
mem[608] = 32'b00111000000000000000000111011111;
mem[609] = 32'b00111111111000000000000000000000;
mem[610] = 32'b00110000000000010000000000000000;
mem[611] = 32'b00110100000000010000000100011011;
mem[612] = 32'b00110000000000010000000000000000;
mem[613] = 32'b00110100000000010000000100011001;
mem[614] = 32'b00110000000000010000000000000000;
mem[615] = 32'b00110100000000010000000100011010;
mem[616] = 32'b00101100000000010000000011010110;
mem[617] = 32'b00001100001001000000000000000000;
mem[618] = 32'b00110000000000010000000000000001;
mem[619] = 32'b00001100001000100000000000000000;
mem[620] = 32'b00001100100000110000000000000000;
mem[621] = 32'b00010000011000100000100000000000;
mem[622] = 32'b00101100001000010000000001001010;
mem[623] = 32'b00110100000000010000000100011100;
mem[624] = 32'b00101100000000010000000011010111;
mem[625] = 32'b00110100000000010000000100011101;
mem[626] = 32'b00110000000000010000000000000000;
mem[627] = 32'b00110100000000010000000100011011;
mem[628] = 32'b00101100000000010000000011111100;
mem[629] = 32'b10011000001000000000000000000000;
mem[630] = 32'b01111100000000010000000000000000;
mem[631] = 32'b00110100000000010000000100011000;
mem[632] = 32'b00101100000000010000000100011011;
mem[633] = 32'b00001100001001000000000000000000;
mem[634] = 32'b00110000000000010000000000000000;
mem[635] = 32'b00001100001001010000000000000000;
mem[636] = 32'b00110000000000010000000000000001;
mem[637] = 32'b00001100001000100000000000000000;
mem[638] = 32'b00001100101000110000000000000000;
mem[639] = 32'b00010000011000100000100000000000;
mem[640] = 32'b00001100001000100000000000000000;
mem[641] = 32'b00001100100000110000000000000000;
mem[642] = 32'b01100000011000100000001010111100;
mem[643] = 32'b00101100000000010000000011111101;
mem[644] = 32'b10011000001000000000000000000000;
mem[645] = 32'b01111100000000010000000000000000;
mem[646] = 32'b00110100000000010000000100011001;
mem[647] = 32'b01111100000000010000000000000000;
mem[648] = 32'b00110100000000010000000100011010;
mem[649] = 32'b00101100000000010000000100011001;
mem[650] = 32'b00001100001101000000000000000000;
mem[651] = 32'b00101100000000010000000100011010;
mem[652] = 32'b00001100001101010000000000000000;
mem[653] = 32'b00101010101101010000010000000000;
mem[654] = 32'b01001010100101010000100000000000;
mem[655] = 32'b00001100001111010000000000000000;
mem[656] = 32'b00110100000000010000000100010111;
mem[657] = 32'b00101100000000010000000100011100;
mem[658] = 32'b00001100001001000000000000000000;
mem[659] = 32'b00101100000000010000000100000111;
mem[660] = 32'b00001100001000100000000000000000;
mem[661] = 32'b00001100100000110000000000000000;
mem[662] = 32'b01011100011000100000001010100001;
mem[663] = 32'b00110000000000010000000000000000;
mem[664] = 32'b00110100000000010000000100011100;
mem[665] = 32'b00101100000000010000000100011101;
mem[666] = 32'b00001100001001000000000000000000;
mem[667] = 32'b00110000000000010000000000000001;
mem[668] = 32'b00001100001000100000000000000000;
mem[669] = 32'b00001100100000110000000000000000;
mem[670] = 32'b00001000011000100000100000000000;
mem[671] = 32'b00110100000000010000000100011101;
mem[672] = 32'b00111000000000000000001010101000;
mem[673] = 32'b00101100000000010000000100011100;
mem[674] = 32'b00001100001001000000000000000000;
mem[675] = 32'b00110000000000010000000000000001;
mem[676] = 32'b00001100001000100000000000000000;
mem[677] = 32'b00001100100000110000000000000000;
mem[678] = 32'b00001000011000100000100000000000;
mem[679] = 32'b00110100000000010000000100011100;
mem[680] = 32'b00101100000000010000000100010111;
mem[681] = 32'b10110100000000010000000000000000;
mem[682] = 32'b00101100000000010000000100011101;
mem[683] = 32'b00001100001000100000000000000000;
mem[684] = 32'b00101100000000010000000100011100;
mem[685] = 32'b00001100001000110000000000000000;
mem[686] = 32'b10011100011000100000000000000000;
mem[687] = 32'b00101100000000010000000100010110;
mem[688] = 32'b00001100001001000000000000000000;
mem[689] = 32'b00110000000000010000000000000001;
mem[690] = 32'b00001100001000100000000000000000;
mem[691] = 32'b00001100100000110000000000000000;
mem[692] = 32'b00001000011000100000100000000000;
mem[693] = 32'b00110100000000010000000100010110;
mem[694] = 32'b10000000000000000000000100010110;
mem[695] = 32'b00101100000000010000000011111110;
mem[696] = 32'b10011000001000000000000000000000;
mem[697] = 32'b01111100000000010000000000000000;
mem[698] = 32'b00110100000000010000000100011011;
mem[699] = 32'b00111000000000000000001001111000;
mem[700] = 32'b00101100000000010000000100010110;
mem[701] = 32'b00001100001001000000000000000000;
mem[702] = 32'b00110000000000010000000000000000;
mem[703] = 32'b00001100001000100000000000000000;
mem[704] = 32'b00001100100000110000000000000000;
mem[705] = 32'b01100000011000100000001011111101;
mem[706] = 32'b00101100000000010000000100000110;
mem[707] = 32'b10011000001000000000000000000000;
mem[708] = 32'b01111100000000010000000000000000;
mem[709] = 32'b00110100000000010000000100011011;
mem[710] = 32'b00101100000000010000000100011011;
mem[711] = 32'b00001100001001000000000000000000;
mem[712] = 32'b00110000000000010000000000000001;
mem[713] = 32'b00001100001000100000000000000000;
mem[714] = 32'b00001100100000110000000000000000;
mem[715] = 32'b01011100011000100000001011111101;
mem[716] = 32'b00101100000000010000000011010110;
mem[717] = 32'b00001100001001000000000000000000;
mem[718] = 32'b00101100000000010000000011010111;
mem[719] = 32'b00110100100000010000000000000100;
mem[720] = 32'b00101100000000010000000011010110;
mem[721] = 32'b00001100001001000000000000000000;
mem[722] = 32'b00101100000000010000000011010110;
mem[723] = 32'b00001100001001010000000000000000;
mem[724] = 32'b00110000000000010000000000000001;
mem[725] = 32'b00001100001000100000000000000000;
mem[726] = 32'b00001100101000110000000000000000;
mem[727] = 32'b00010000011000100000100000000000;
mem[728] = 32'b00101100001000010000000001001010;
mem[729] = 32'b00001100001001010000000000000000;
mem[730] = 32'b00110000000000010000000000000001;
mem[731] = 32'b00001100001000100000000000000000;
mem[732] = 32'b00001100101000110000000000000000;
mem[733] = 32'b00001000011000100000100000000000;
mem[734] = 32'b00110100100000010000000000100111;
mem[735] = 32'b00101100000000010000000011010110;
mem[736] = 32'b00001100001001000000000000000000;
mem[737] = 32'b00101100000000010000000100011100;
mem[738] = 32'b00001100001001010000000000000000;
mem[739] = 32'b00110000000000010000000000000001;
mem[740] = 32'b00001100001000100000000000000000;
mem[741] = 32'b00001100101000110000000000000000;
mem[742] = 32'b00010000011000100000100000000000;
mem[743] = 32'b00110100100000010000000001001010;
mem[744] = 32'b00101100000000010000000011010110;
mem[745] = 32'b00001100001001000000000000000000;
mem[746] = 32'b00101100000000010000000100011000;
mem[747] = 32'b00110100100000010000000001101101;
mem[748] = 32'b00101100000000010000000011010110;
mem[749] = 32'b00001100001001000000000000000000;
mem[750] = 32'b00110000000000010000000000000001;
mem[751] = 32'b00110100100000010000000010010000;
mem[752] = 32'b00101100000000010000000011010110;
mem[753] = 32'b00001100001001000000000000000000;
mem[754] = 32'b00101100000000010000000100010110;
mem[755] = 32'b00110100100000010000000010110011;
mem[756] = 32'b00101100000000010000000011010110;
mem[757] = 32'b00001100001001000000000000000000;
mem[758] = 32'b00110000000000010000000000000001;
mem[759] = 32'b00001100001000100000000000000000;
mem[760] = 32'b00001100100000110000000000000000;
mem[761] = 32'b00001000011000100000100000000000;
mem[762] = 32'b00110100000000010000000011010110;
mem[763] = 32'b00101100000000010000000100011101;
mem[764] = 32'b00110100000000010000000011010111;
mem[765] = 32'b00111111111000000000000000000000;
mem[766] = 32'b00110000000000010000000000000100;
mem[767] = 32'b00110100000000010000000100011110;
mem[768] = 32'b00101100000000010000000100011110;
mem[769] = 32'b10110100000000010000000000000000;
mem[770] = 32'b00111111111000000000000000000000;
mem[771] = 32'b10110000000000010000000000000000;
mem[772] = 32'b00110100000000010000000100011111;
mem[773] = 32'b10000000000000000000000100011111;
mem[774] = 32'b00111111111000000000000000000000;
mem[775] = 32'b00001111110111101111111111111111;
mem[776] = 32'b00110111110111110000000000000000;
mem[777] = 32'b00101100000000010000000100100000;
mem[778] = 32'b00110100000000010000000101011011;
mem[779] = 32'b00101100000000010000000101011011;
mem[780] = 32'b00110100000000010000000100001101;
mem[781] = 32'b10000100000000000000000110000010;
mem[782] = 32'b00101111110111110000000000000000;
mem[783] = 32'b00001111110111100000000000000001;
mem[784] = 32'b00001111101000010000000000000000;
mem[785] = 32'b00110100000000010000000100100001;
mem[786] = 32'b00101100000000010000000100100001;
mem[787] = 32'b00001100001001000000000000000000;
mem[788] = 32'b00110000000000010000000000000000;
mem[789] = 32'b00001100001000100000000000000000;
mem[790] = 32'b00001100100000110000000000000000;
mem[791] = 32'b01100000011000100000001101001111;
mem[792] = 32'b00110000000000010000000000000000;
mem[793] = 32'b00110100000000010000000100100100;
mem[794] = 32'b00101100000000010000000100100001;
mem[795] = 32'b00101100001000010000000000100111;
mem[796] = 32'b00110100000000010000000100100010;
mem[797] = 32'b00101100000000010000000100100001;
mem[798] = 32'b00101100001000010000000000000100;
mem[799] = 32'b00110100000000010000000100100011;
mem[800] = 32'b00000000000000000000000000000000;
mem[801] = 32'b00101100000000010000000100100100;
mem[802] = 32'b00001100001001000000000000000000;
mem[803] = 32'b00101100000000010000000100100001;
mem[804] = 32'b00101100001000010000000010110011;
mem[805] = 32'b00001100001000100000000000000000;
mem[806] = 32'b00001100100000110000000000000000;
mem[807] = 32'b01110000011000100000001101001111;
mem[808] = 32'b00101100000000010000000100100011;
mem[809] = 32'b00001100001000100000000000000000;
mem[810] = 32'b00101100000000010000000100100010;
mem[811] = 32'b00001100001000110000000000000000;
mem[812] = 32'b00110000000000010000000000000001;
mem[813] = 32'b10010100000000010000000000000000;
mem[814] = 32'b10001000011000100000000000000000;
mem[815] = 32'b10010100000000000000000000000000;
mem[816] = 32'b00101100000000010000000100100010;
mem[817] = 32'b00001100001001000000000000000000;
mem[818] = 32'b00101100000000010000000100000111;
mem[819] = 32'b00001100001000100000000000000000;
mem[820] = 32'b00001100100000110000000000000000;
mem[821] = 32'b01011100011000100000001101000000;
mem[822] = 32'b00110000000000010000000000000000;
mem[823] = 32'b00110100000000010000000100100010;
mem[824] = 32'b00101100000000010000000100100011;
mem[825] = 32'b00001100001001000000000000000000;
mem[826] = 32'b00110000000000010000000000000001;
mem[827] = 32'b00001100001000100000000000000000;
mem[828] = 32'b00001100100000110000000000000000;
mem[829] = 32'b00001000011000100000100000000000;
mem[830] = 32'b00110100000000010000000100100011;
mem[831] = 32'b00111000000000000000001101000111;
mem[832] = 32'b00101100000000010000000100100010;
mem[833] = 32'b00001100001001000000000000000000;
mem[834] = 32'b00110000000000010000000000000001;
mem[835] = 32'b00001100001000100000000000000000;
mem[836] = 32'b00001100100000110000000000000000;
mem[837] = 32'b00001000011000100000100000000000;
mem[838] = 32'b00110100000000010000000100100010;
mem[839] = 32'b00101100000000010000000100100100;
mem[840] = 32'b00001100001001000000000000000000;
mem[841] = 32'b00110000000000010000000000000001;
mem[842] = 32'b00001100001000100000000000000000;
mem[843] = 32'b00001100100000110000000000000000;
mem[844] = 32'b00001000011000100000100000000000;
mem[845] = 32'b00110100000000010000000100100100;
mem[846] = 32'b00111000000000000000001100100001;
mem[847] = 32'b00111111111000000000000000000000;
mem[848] = 32'b00101100000000010000000100100101;
mem[849] = 32'b00001100001110100000000000000000;
mem[850] = 32'b00110000000110110000000000100000;
mem[851] = 32'b00011011010110111101100000000000;
mem[852] = 32'b00001111010110100000000000000001;
mem[853] = 32'b11000111011000010000000101011110;
mem[854] = 32'b00001111011110110000000000000001;
mem[855] = 32'b11000111011000100000000101011110;
mem[856] = 32'b00001111011110110000000000000001;
mem[857] = 32'b11000111011000110000000101011110;
mem[858] = 32'b00001111011110110000000000000001;
mem[859] = 32'b11000111011001000000000101011110;
mem[860] = 32'b00001111011110110000000000000001;
mem[861] = 32'b11000111011001010000000101011110;
mem[862] = 32'b00001111011110110000000000000001;
mem[863] = 32'b11000111011111010000000101011110;
mem[864] = 32'b00001111011110110000000000000001;
mem[865] = 32'b11000111011111100000000101011110;
mem[866] = 32'b00001111011110110000000000000001;
mem[867] = 32'b11000111011111110000000101011110;
mem[868] = 32'b00001111011110110000000000000001;
mem[869] = 32'b00111111111000000000000000000000;
mem[870] = 32'b00101100000000010000000100100110;
mem[871] = 32'b00001100001110100000000000000000;
mem[872] = 32'b00110000000110110000000000100000;
mem[873] = 32'b00011011010110111101100000000000;
mem[874] = 32'b00001111010110100000000000000001;
mem[875] = 32'b11001011011000010000000101011110;
mem[876] = 32'b00001111011110110000000000000001;
mem[877] = 32'b11001011011000100000000101011110;
mem[878] = 32'b00001111011110110000000000000001;
mem[879] = 32'b11001011011000110000000101011110;
mem[880] = 32'b00001111011110110000000000000001;
mem[881] = 32'b11001011011001000000000101011110;
mem[882] = 32'b00001111011110110000000000000001;
mem[883] = 32'b11001011011001010000000101011110;
mem[884] = 32'b00001111011110110000000000000001;
mem[885] = 32'b11001011011111010000000101011110;
mem[886] = 32'b00001111011110110000000000000001;
mem[887] = 32'b11001011011111100000000101011110;
mem[888] = 32'b00001111011110110000000000000001;
mem[889] = 32'b11001011011111110000000101011110;
mem[890] = 32'b00001111011110110000000000000001;
mem[891] = 32'b00111111111000000000000000000000;
mem[892] = 32'b00110000000000010000000000000000;
mem[893] = 32'b00110100000000010000000100101000;
mem[894] = 32'b00110000000000010000000000000100;
mem[895] = 32'b00110100000000010000000100001001;
mem[896] = 32'b00101100000000010000000100101000;
mem[897] = 32'b00001100001001000000000000000000;
mem[898] = 32'b00110000000000010000000000110010;
mem[899] = 32'b00110100100000010000000011011001;
mem[900] = 32'b00101100000000010000000100101000;
mem[901] = 32'b00001100001001000000000000000000;
mem[902] = 32'b00101100000000010000000100101000;
mem[903] = 32'b00001100001001010000000000000000;
mem[904] = 32'b00110000000000010000000000000001;
mem[905] = 32'b00001100001000100000000000000000;
mem[906] = 32'b00001100101000110000000000000000;
mem[907] = 32'b00001000011000100000100000000000;
mem[908] = 32'b00110100100000010000000011100011;
mem[909] = 32'b00101100000000010000000100101000;
mem[910] = 32'b00001100001001000000000000000000;
mem[911] = 32'b00110000000000010000000000000000;
mem[912] = 32'b00110100100000010000000011101101;
mem[913] = 32'b00101100000000010000000100101000;
mem[914] = 32'b00001100001001000000000000000000;
mem[915] = 32'b00110000000000010000000000000001;
mem[916] = 32'b00001100001000100000000000000000;
mem[917] = 32'b00001100100000110000000000000000;
mem[918] = 32'b00001000011000100000100000000000;
mem[919] = 32'b00110100000000010000000100101000;
mem[920] = 32'b00101100000000010000000100101000;
mem[921] = 32'b00001100001001000000000000000000;
mem[922] = 32'b00110000000000010000000000110011;
mem[923] = 32'b00110100100000010000000011011001;
mem[924] = 32'b00101100000000010000000100101000;
mem[925] = 32'b00001100001001000000000000000000;
mem[926] = 32'b00101100000000010000000100101000;
mem[927] = 32'b00001100001001010000000000000000;
mem[928] = 32'b00110000000000010000000000000001;
mem[929] = 32'b00001100001000100000000000000000;
mem[930] = 32'b00001100101000110000000000000000;
mem[931] = 32'b00001000011000100000100000000000;
mem[932] = 32'b00110100100000010000000011100011;
mem[933] = 32'b00101100000000010000000100101000;
mem[934] = 32'b00001100001001000000000000000000;
mem[935] = 32'b00110000000000010000000000000000;
mem[936] = 32'b00110100100000010000000011101101;
mem[937] = 32'b00101100000000010000000100101000;
mem[938] = 32'b00001100001001000000000000000000;
mem[939] = 32'b00110000000000010000000000000001;
mem[940] = 32'b00001100001000100000000000000000;
mem[941] = 32'b00001100100000110000000000000000;
mem[942] = 32'b00001000011000100000100000000000;
mem[943] = 32'b00110100000000010000000100101000;
mem[944] = 32'b00101100000000010000000100101000;
mem[945] = 32'b00001100001001000000000000000000;
mem[946] = 32'b00110000000000010000000000110100;
mem[947] = 32'b00110100100000010000000011011001;
mem[948] = 32'b00101100000000010000000100101000;
mem[949] = 32'b00001100001001000000000000000000;
mem[950] = 32'b00101100000000010000000100101000;
mem[951] = 32'b00001100001001010000000000000000;
mem[952] = 32'b00110000000000010000000000000001;
mem[953] = 32'b00001100001000100000000000000000;
mem[954] = 32'b00001100101000110000000000000000;
mem[955] = 32'b00001000011000100000100000000000;
mem[956] = 32'b00110100100000010000000011100011;
mem[957] = 32'b00101100000000010000000100101000;
mem[958] = 32'b00001100001001000000000000000000;
mem[959] = 32'b00110000000000010000000000000000;
mem[960] = 32'b00110100100000010000000011101101;
mem[961] = 32'b00101100000000010000000100101000;
mem[962] = 32'b00001100001001000000000000000000;
mem[963] = 32'b00110000000000010000000000000001;
mem[964] = 32'b00001100001000100000000000000000;
mem[965] = 32'b00001100100000110000000000000000;
mem[966] = 32'b00001000011000100000100000000000;
mem[967] = 32'b00110100000000010000000100101000;
mem[968] = 32'b00101100000000010000000100101000;
mem[969] = 32'b00001100001001000000000000000000;
mem[970] = 32'b00110000000000010000000000110101;
mem[971] = 32'b00110100100000010000000011011001;
mem[972] = 32'b00101100000000010000000100101000;
mem[973] = 32'b00001100001001000000000000000000;
mem[974] = 32'b00101100000000010000000100101000;
mem[975] = 32'b00001100001001010000000000000000;
mem[976] = 32'b00110000000000010000000000000001;
mem[977] = 32'b00001100001000100000000000000000;
mem[978] = 32'b00001100101000110000000000000000;
mem[979] = 32'b00001000011000100000100000000000;
mem[980] = 32'b00110100100000010000000011100011;
mem[981] = 32'b00101100000000010000000100101000;
mem[982] = 32'b00001100001001000000000000000000;
mem[983] = 32'b00110000000000010000000000000000;
mem[984] = 32'b00110100100000010000000011101101;
mem[985] = 32'b00101100000000010000000100101000;
mem[986] = 32'b00001100001001000000000000000000;
mem[987] = 32'b00110000000000010000000000000001;
mem[988] = 32'b00001100001000100000000000000000;
mem[989] = 32'b00001100100000110000000000000000;
mem[990] = 32'b00001000011000100000100000000000;
mem[991] = 32'b00110100000000010000000100101000;
mem[992] = 32'b00101100000000010000000100101000;
mem[993] = 32'b00001100001001000000000000000000;
mem[994] = 32'b00110000000000010000000000001010;
mem[995] = 32'b00001100001000100000000000000000;
mem[996] = 32'b00001100100000110000000000000000;
mem[997] = 32'b01110000011000100000001111111010;
mem[998] = 32'b00101100000000010000000100101000;
mem[999] = 32'b00001100001001000000000000000000;
mem[1000] = 32'b00110000000000010000000000000000;
mem[1001] = 32'b00110100100000010000000011011001;
mem[1002] = 32'b00101100000000010000000100101000;
mem[1003] = 32'b00001100001001000000000000000000;
mem[1004] = 32'b00110000000000010000000000000000;
mem[1005] = 32'b00110100100000010000000011100011;
mem[1006] = 32'b00101100000000010000000100101000;
mem[1007] = 32'b00001100001001000000000000000000;
mem[1008] = 32'b00110000000000010000000000000000;
mem[1009] = 32'b00110100100000010000000011101101;
mem[1010] = 32'b00101100000000010000000100101000;
mem[1011] = 32'b00001100001001000000000000000000;
mem[1012] = 32'b00110000000000010000000000000001;
mem[1013] = 32'b00001100001000100000000000000000;
mem[1014] = 32'b00001100100000110000000000000000;
mem[1015] = 32'b00001000011000100000100000000000;
mem[1016] = 32'b00110100000000010000000100101000;
mem[1017] = 32'b00111000000000000000001111100000;
mem[1018] = 32'b00111111111000000000000000000000;
mem[1019] = 32'b00110000000000010000000000000000;
mem[1020] = 32'b00110100000000010000000100101001;
mem[1021] = 32'b00110000000000010000000000000001;
mem[1022] = 32'b00110100000000010000000100101100;
mem[1023] = 32'b00110000000000010000000000000000;
mem[1024] = 32'b00110100000000010000000100101110;
mem[1025] = 32'b00001111110111101111111111111111;
mem[1026] = 32'b00110111110111110000000000000000;
mem[1027] = 32'b10000100000000000000001101111100;
mem[1028] = 32'b00101111110111110000000000000000;
mem[1029] = 32'b00001111110111100000000000000001;
mem[1030] = 32'b00110000000000010000000000101000;
mem[1031] = 32'b10111100000000010000000000000000;
mem[1032] = 32'b00101100000000010000000100001001;
mem[1033] = 32'b00110100000000010000000100101011;
mem[1034] = 32'b00110000000000010000000000000000;
mem[1035] = 32'b10100100001000000000000000000000;
mem[1036] = 32'b00101100000000010000000100101011;
mem[1037] = 32'b00001100001001000000000000000000;
mem[1038] = 32'b00110000000000010000000000000000;
mem[1039] = 32'b00001100001000100000000000000000;
mem[1040] = 32'b00001100100000110000000000000000;
mem[1041] = 32'b01101100011000100000010100011011;
mem[1042] = 32'b00101100000000010000000100101100;
mem[1043] = 32'b00001100001001000000000000000000;
mem[1044] = 32'b00110000000000010000000000000000;
mem[1045] = 32'b00001100001000100000000000000000;
mem[1046] = 32'b00001100100000110000000000000000;
mem[1047] = 32'b01100000011000100000010010101011;
mem[1048] = 32'b00101100000000010000000100101110;
mem[1049] = 32'b00001100001001000000000000000000;
mem[1050] = 32'b00110000000000010000000000000001;
mem[1051] = 32'b00001100001000100000000000000000;
mem[1052] = 32'b00001100100000110000000000000000;
mem[1053] = 32'b01011100011000100000010001110001;
mem[1054] = 32'b00101100000000010000000100101001;
mem[1055] = 32'b00001100001001000000000000000000;
mem[1056] = 32'b00101100000000010000000100101011;
mem[1057] = 32'b00001100001001010000000000000000;
mem[1058] = 32'b00110000000000010000000000000001;
mem[1059] = 32'b00001100001000100000000000000000;
mem[1060] = 32'b00001100101000110000000000000000;
mem[1061] = 32'b00010000011000100000100000000000;
mem[1062] = 32'b00001100001000100000000000000000;
mem[1063] = 32'b00001100100000110000000000000000;
mem[1064] = 32'b01110000011000100000010001011100;
mem[1065] = 32'b00101100000000010000000100101001;
mem[1066] = 32'b00110100000000010000000100101101;
mem[1067] = 32'b00101100000000010000000100101101;
mem[1068] = 32'b00001100001001000000000000000000;
mem[1069] = 32'b00101100000000010000000100101011;
mem[1070] = 32'b00001100001001010000000000000000;
mem[1071] = 32'b00110000000000010000000000000001;
mem[1072] = 32'b00001100001000100000000000000000;
mem[1073] = 32'b00001100101000110000000000000000;
mem[1074] = 32'b00010000011000100000100000000000;
mem[1075] = 32'b00001100001000100000000000000000;
mem[1076] = 32'b00001100100000110000000000000000;
mem[1077] = 32'b01110000011000100000010001011100;
mem[1078] = 32'b00101100000000010000000100101101;
mem[1079] = 32'b00001100001001000000000000000000;
mem[1080] = 32'b00101100000000010000000100101101;
mem[1081] = 32'b00001100001001010000000000000000;
mem[1082] = 32'b00110000000000010000000000000001;
mem[1083] = 32'b00001100001000100000000000000000;
mem[1084] = 32'b00001100101000110000000000000000;
mem[1085] = 32'b00001000011000100000100000000000;
mem[1086] = 32'b00101100001000010000000011101101;
mem[1087] = 32'b00110100100000010000000011101101;
mem[1088] = 32'b00101100000000010000000100101101;
mem[1089] = 32'b00001100001001000000000000000000;
mem[1090] = 32'b00101100000000010000000100101101;
mem[1091] = 32'b00001100001001010000000000000000;
mem[1092] = 32'b00110000000000010000000000000001;
mem[1093] = 32'b00001100001000100000000000000000;
mem[1094] = 32'b00001100101000110000000000000000;
mem[1095] = 32'b00001000011000100000100000000000;
mem[1096] = 32'b00101100001000010000000011011001;
mem[1097] = 32'b00110100100000010000000011011001;
mem[1098] = 32'b00101100000000010000000100101101;
mem[1099] = 32'b00001100001001000000000000000000;
mem[1100] = 32'b00101100000000010000000100101101;
mem[1101] = 32'b00001100001001010000000000000000;
mem[1102] = 32'b00110000000000010000000000000001;
mem[1103] = 32'b00001100001000100000000000000000;
mem[1104] = 32'b00001100101000110000000000000000;
mem[1105] = 32'b00001000011000100000100000000000;
mem[1106] = 32'b00101100001000010000000011100011;
mem[1107] = 32'b00110100100000010000000011100011;
mem[1108] = 32'b00101100000000010000000100101101;
mem[1109] = 32'b00001100001001000000000000000000;
mem[1110] = 32'b00110000000000010000000000000001;
mem[1111] = 32'b00001100001000100000000000000000;
mem[1112] = 32'b00001100100000110000000000000000;
mem[1113] = 32'b00001000011000100000100000000000;
mem[1114] = 32'b00110100000000010000000100101101;
mem[1115] = 32'b00111000000000000000010000101011;
mem[1116] = 32'b00101100000000010000000100101001;
mem[1117] = 32'b00001100001001000000000000000000;
mem[1118] = 32'b00101100000000010000000100101011;
mem[1119] = 32'b00001100001001010000000000000000;
mem[1120] = 32'b00110000000000010000000000000001;
mem[1121] = 32'b00001100001000100000000000000000;
mem[1122] = 32'b00001100101000110000000000000000;
mem[1123] = 32'b00010000011000100000100000000000;
mem[1124] = 32'b00001100001000100000000000000000;
mem[1125] = 32'b00001100100000110000000000000000;
mem[1126] = 32'b01011100011000100000010001101001;
mem[1127] = 32'b00110000000000010000000000000000;
mem[1128] = 32'b00110100000000010000000100101001;
mem[1129] = 32'b00101100000000010000000100101011;
mem[1130] = 32'b00001100001001000000000000000000;
mem[1131] = 32'b00110000000000010000000000000001;
mem[1132] = 32'b00001100001000100000000000000000;
mem[1133] = 32'b00001100100000110000000000000000;
mem[1134] = 32'b00010000011000100000100000000000;
mem[1135] = 32'b00110100000000010000000100101011;
mem[1136] = 32'b00111000000000000000010010011001;
mem[1137] = 32'b00101100000000010000000100101001;
mem[1138] = 32'b00001100001001000000000000000000;
mem[1139] = 32'b00110000000000010000000000000000;
mem[1140] = 32'b00001100001000100000000000000000;
mem[1141] = 32'b00001100100000110000000000000000;
mem[1142] = 32'b01011100011000100000010001111111;
mem[1143] = 32'b00101100000000010000000100101011;
mem[1144] = 32'b00001100001001000000000000000000;
mem[1145] = 32'b00110000000000010000000000000001;
mem[1146] = 32'b00001100001000100000000000000000;
mem[1147] = 32'b00001100100000110000000000000000;
mem[1148] = 32'b00010000011000100000100000000000;
mem[1149] = 32'b00110100000000010000000100101111;
mem[1150] = 32'b00111000000000000000010010000110;
mem[1151] = 32'b00101100000000010000000100101001;
mem[1152] = 32'b00001100001001000000000000000000;
mem[1153] = 32'b00110000000000010000000000000001;
mem[1154] = 32'b00001100001000100000000000000000;
mem[1155] = 32'b00001100100000110000000000000000;
mem[1156] = 32'b00010000011000100000100000000000;
mem[1157] = 32'b00110100000000010000000100101111;
mem[1158] = 32'b00101100000000010000000100101111;
mem[1159] = 32'b00001100001001000000000000000000;
mem[1160] = 32'b10100000000000010000000000000000;
mem[1161] = 32'b00110100100000010000000011101101;
mem[1162] = 32'b00001111110111101111111111111111;
mem[1163] = 32'b00110111110111110000000000000000;
mem[1164] = 32'b00101100000000010000000100101111;
mem[1165] = 32'b00101100001000010000000011100011;
mem[1166] = 32'b00001100001001000000000000000000;
mem[1167] = 32'b00110000000000010000000000000001;
mem[1168] = 32'b00001100001000100000000000000000;
mem[1169] = 32'b00001100100000110000000000000000;
mem[1170] = 32'b00010000011000100000100000000000;
mem[1171] = 32'b00110100000000010000000101011011;
mem[1172] = 32'b00101100000000010000000101011011;
mem[1173] = 32'b00110100000000010000000100100110;
mem[1174] = 32'b10000100000000000000001101100110;
mem[1175] = 32'b00101111110111110000000000000000;
mem[1176] = 32'b00001111110111100000000000000001;
mem[1177] = 32'b00001111110111101111111111111111;
mem[1178] = 32'b00110111110111110000000000000000;
mem[1179] = 32'b00101100000000010000000100101001;
mem[1180] = 32'b00101100001000010000000011100011;
mem[1181] = 32'b00001100001001000000000000000000;
mem[1182] = 32'b00110000000000010000000000000001;
mem[1183] = 32'b00001100001000100000000000000000;
mem[1184] = 32'b00001100100000110000000000000000;
mem[1185] = 32'b00010000011000100000100000000000;
mem[1186] = 32'b00110100000000010000000101011011;
mem[1187] = 32'b00101100000000010000000101011011;
mem[1188] = 32'b00110100000000010000000100100101;
mem[1189] = 32'b10000100000000000000001101010000;
mem[1190] = 32'b00101111110111110000000000000000;
mem[1191] = 32'b00001111110111100000000000000001;
mem[1192] = 32'b00101100000000010000000100101001;
mem[1193] = 32'b00101100001000010000000011101101;
mem[1194] = 32'b10100100001000000000000000000000;
mem[1195] = 32'b00101100000000010000000100101001;
mem[1196] = 32'b00101100001000010000000011100011;
mem[1197] = 32'b00110100000000010000000100110000;
mem[1198] = 32'b00101100000000010000000000000010;
mem[1199] = 32'b00001100001001000000000000000000;
mem[1200] = 32'b00110000000000010000000000000000;
mem[1201] = 32'b00001100001000100000000000000000;
mem[1202] = 32'b00001100100000110000000000000000;
mem[1203] = 32'b01011100011000100000010010110101;
mem[1204] = 32'b11000000000000000000000000000000;
mem[1205] = 32'b00101100000000010000000000000010;
mem[1206] = 32'b00001100001001000000000000000000;
mem[1207] = 32'b00110000000000010000000000000011;
mem[1208] = 32'b00001100001000100000000000000000;
mem[1209] = 32'b00001100100000110000000000000000;
mem[1210] = 32'b01011100011000100000010010111100;
mem[1211] = 32'b11000000000000000000000000000000;
mem[1212] = 32'b00101100000100110000000100110000;
mem[1213] = 32'b10010100000100110000000000000000;
mem[1214] = 32'b00101100000100110000000100110000;
mem[1215] = 32'b10001100000100110000000000000000;
mem[1216] = 32'b10101100000000000000000000000000;
mem[1217] = 32'b00000000000000000000000000000000;
mem[1218] = 32'b00110000000100110000000000000000;
mem[1219] = 32'b10010100000100110000000000000000;
mem[1220] = 32'b00110000000100110000000000000000;
mem[1221] = 32'b10001100000100110000000000000000;
mem[1222] = 32'b10101000000000000000100000000000;
mem[1223] = 32'b00110100000000010000000000000010;
mem[1224] = 32'b00101100000000010000000000000010;
mem[1225] = 32'b00001100001001000000000000000000;
mem[1226] = 32'b00110000000000010000000000000000;
mem[1227] = 32'b00001100001000100000000000000000;
mem[1228] = 32'b00001100100000110000000000000000;
mem[1229] = 32'b01011100011000100000010011101000;
mem[1230] = 32'b00110000000000010000000000000000;
mem[1231] = 32'b00110100000000010000000100101110;
mem[1232] = 32'b00110000000000010000000000000001;
mem[1233] = 32'b00110100000000010000000100101100;
mem[1234] = 32'b00101100000000010000000100101001;
mem[1235] = 32'b00001100001001000000000000000000;
mem[1236] = 32'b00101100000000010000000100101011;
mem[1237] = 32'b00001100001001010000000000000000;
mem[1238] = 32'b00110000000000010000000000000001;
mem[1239] = 32'b00001100001000100000000000000000;
mem[1240] = 32'b00001100101000110000000000000000;
mem[1241] = 32'b00010000011000100000100000000000;
mem[1242] = 32'b00001100001000100000000000000000;
mem[1243] = 32'b00001100100000110000000000000000;
mem[1244] = 32'b01011100011000100000010011100000;
mem[1245] = 32'b00110000000000010000000000000000;
mem[1246] = 32'b00110100000000010000000100101001;
mem[1247] = 32'b00111000000000000000010011100111;
mem[1248] = 32'b00101100000000010000000100101001;
mem[1249] = 32'b00001100001001000000000000000000;
mem[1250] = 32'b00110000000000010000000000000001;
mem[1251] = 32'b00001100001000100000000000000000;
mem[1252] = 32'b00001100100000110000000000000000;
mem[1253] = 32'b00001000011000100000100000000000;
mem[1254] = 32'b00110100000000010000000100101001;
mem[1255] = 32'b00111000000000000000010100011010;
mem[1256] = 32'b00101100000000010000000000000010;
mem[1257] = 32'b00001100001001000000000000000000;
mem[1258] = 32'b00110000000000010000000000000001;
mem[1259] = 32'b00001100001000100000000000000000;
mem[1260] = 32'b00001100100000110000000000000000;
mem[1261] = 32'b01011100011000100000010011111000;
mem[1262] = 32'b00110000000000010000000000000000;
mem[1263] = 32'b00110100000000010000000100101110;
mem[1264] = 32'b00110000000000010000000000000000;
mem[1265] = 32'b00110100000000010000000100101100;
mem[1266] = 32'b00001111110111101111111111111111;
mem[1267] = 32'b00110111110111110000000000000000;
mem[1268] = 32'b10000100000000000000001011111110;
mem[1269] = 32'b00101111110111110000000000000000;
mem[1270] = 32'b00001111110111100000000000000001;
mem[1271] = 32'b00111000000000000000010100011010;
mem[1272] = 32'b00101100000000010000000000000010;
mem[1273] = 32'b00001100001001000000000000000000;
mem[1274] = 32'b00110000000000010000000000000010;
mem[1275] = 32'b00001100001000100000000000000000;
mem[1276] = 32'b00001100100000110000000000000000;
mem[1277] = 32'b01011100011000100000010100001000;
mem[1278] = 32'b00110000000000010000000000000000;
mem[1279] = 32'b00110100000000010000000100101110;
mem[1280] = 32'b00110000000000010000000000000000;
mem[1281] = 32'b00110100000000010000000100101100;
mem[1282] = 32'b00001111110111101111111111111111;
mem[1283] = 32'b00110111110111110000000000000000;
mem[1284] = 32'b10000100000000000000001100000011;
mem[1285] = 32'b00101111110111110000000000000000;
mem[1286] = 32'b00001111110111100000000000000001;
mem[1287] = 32'b00111000000000000000010100011010;
mem[1288] = 32'b00101100000000010000000000000010;
mem[1289] = 32'b00001100001001000000000000000000;
mem[1290] = 32'b00110000000000010000000000000011;
mem[1291] = 32'b00001100001000100000000000000000;
mem[1292] = 32'b00001100100000110000000000000000;
mem[1293] = 32'b01011100011000100000010100011010;
mem[1294] = 32'b00110000000000010000000000000001;
mem[1295] = 32'b00110100000000010000000100101110;
mem[1296] = 32'b00110000000000010000000000000001;
mem[1297] = 32'b00110100000000010000000100101100;
mem[1298] = 32'b00101100000000010000000100101011;
mem[1299] = 32'b00001100001001000000000000000000;
mem[1300] = 32'b00110000000000010000000000000001;
mem[1301] = 32'b00001100001000100000000000000000;
mem[1302] = 32'b00001100100000110000000000000000;
mem[1303] = 32'b01011100011000100000010100011010;
mem[1304] = 32'b00110000000000010000000000000000;
mem[1305] = 32'b00110100000000010000000100101011;
mem[1306] = 32'b00111000000000000000010000001100;
mem[1307] = 32'b00111111111000000000000000000000;
mem[1308] = 32'b00110000000000010000000000001010;
mem[1309] = 32'b00110100000000010000000100110001;
mem[1310] = 32'b10000100000000000000001111111011;
mem[1311] = 32'b00000100000000000000000000000000;

mem[1*(ADDR_WIDTH)+0] =  32'b00000000000000000000000000000000;
mem[1*(ADDR_WIDTH)+1] =  32'b00111000000000000000000000100110;
mem[1*(ADDR_WIDTH)+2] =  32'b00110000000000010000000000000000;
mem[1*(ADDR_WIDTH)+3] =  32'b00110100000000010000000000010110;
mem[1*(ADDR_WIDTH)+4] =  32'b00110000000000010000000000000000;
mem[1*(ADDR_WIDTH)+5] =  32'b00110100000000010000000000010111;
mem[1*(ADDR_WIDTH)+6] =  32'b00101100000000010000000000010111;
mem[1*(ADDR_WIDTH)+7] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+8] =  32'b00101100000000010000000000010101;
mem[1*(ADDR_WIDTH)+9] =  32'b00001100001000100000000000000000;
mem[1*(ADDR_WIDTH)+10] =  32'b00001100100000110000000000000000;
mem[1*(ADDR_WIDTH)+11] =  32'b01110000011000100000000000011110;
mem[1*(ADDR_WIDTH)+12] =  32'b00101100000000010000000000010110;
mem[1*(ADDR_WIDTH)+13] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+14] =  32'b00101100000000010000000000010111;
mem[1*(ADDR_WIDTH)+15] =  32'b00101100000000100000000000010100;
mem[1*(ADDR_WIDTH)+16] =  32'b00001000010000010000100000000000;
mem[1*(ADDR_WIDTH)+17] =  32'b00101100001000010000000000000000;
mem[1*(ADDR_WIDTH)+18] =  32'b00001100001000100000000000000000;
mem[1*(ADDR_WIDTH)+19] =  32'b00001100100000110000000000000000;
mem[1*(ADDR_WIDTH)+20] =  32'b00001000011000100000100000000000;
mem[1*(ADDR_WIDTH)+21] =  32'b00110100000000010000000000010110;
mem[1*(ADDR_WIDTH)+22] =  32'b00101100000000010000000000010111;
mem[1*(ADDR_WIDTH)+23] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+24] =  32'b00110000000000010000000000000001;
mem[1*(ADDR_WIDTH)+25] =  32'b00001100001000100000000000000000;
mem[1*(ADDR_WIDTH)+26] =  32'b00001100100000110000000000000000;
mem[1*(ADDR_WIDTH)+27] =  32'b00001000011000100000100000000000;
mem[1*(ADDR_WIDTH)+28] =  32'b00110100000000010000000000010111;
mem[1*(ADDR_WIDTH)+29] =  32'b00111000000000000000000000000110;
mem[1*(ADDR_WIDTH)+30] =  32'b00101100000000010000000000010110;
mem[1*(ADDR_WIDTH)+31] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+32] =  32'b00101100000000010000000000010101;
mem[1*(ADDR_WIDTH)+33] =  32'b00001100001000100000000000000000;
mem[1*(ADDR_WIDTH)+34] =  32'b00001100100000110000000000000000;
mem[1*(ADDR_WIDTH)+35] =  32'b00011100011000100000100000000000;
mem[1*(ADDR_WIDTH)+36] =  32'b00001100001111010000000000000000;
mem[1*(ADDR_WIDTH)+37] =  32'b00111111111000000000000000000000;
mem[1*(ADDR_WIDTH)+38] =  32'b00110000000000010000000000000000;
mem[1*(ADDR_WIDTH)+39] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+40] =  32'b00110000000000010000000000000101;
mem[1*(ADDR_WIDTH)+41] =  32'b00110100100000010000000000000000;
mem[1*(ADDR_WIDTH)+42] =  32'b00110000000000010000000000000001;
mem[1*(ADDR_WIDTH)+43] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+44] =  32'b00110000000000010000000000000111;
mem[1*(ADDR_WIDTH)+45] =  32'b00110100100000010000000000000000;
mem[1*(ADDR_WIDTH)+46] =  32'b00110000000000010000000000000010;
mem[1*(ADDR_WIDTH)+47] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+48] =  32'b00110000000000010000000000000010;
mem[1*(ADDR_WIDTH)+49] =  32'b00110100100000010000000000000000;
mem[1*(ADDR_WIDTH)+50] =  32'b00110000000000010000000000000011;
mem[1*(ADDR_WIDTH)+51] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+52] =  32'b00110000000000010000000000001100;
mem[1*(ADDR_WIDTH)+53] =  32'b00110100100000010000000000000000;
mem[1*(ADDR_WIDTH)+54] =  32'b00110000000000010000000000000100;
mem[1*(ADDR_WIDTH)+55] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+56] =  32'b00110000000000010000000000010010;
mem[1*(ADDR_WIDTH)+57] =  32'b00110100100000010000000000000000;
mem[1*(ADDR_WIDTH)+58] =  32'b00110000000000010000000000000101;
mem[1*(ADDR_WIDTH)+59] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+60] =  32'b00110000000000010000000000000001;
mem[1*(ADDR_WIDTH)+61] =  32'b00110100100000010000000000000000;
mem[1*(ADDR_WIDTH)+62] =  32'b00110000000000010000000000000110;
mem[1*(ADDR_WIDTH)+63] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+64] =  32'b00110000000000010000000000000010;
mem[1*(ADDR_WIDTH)+65] =  32'b00110100100000010000000000000000;
mem[1*(ADDR_WIDTH)+66] =  32'b00110000000000010000000000000111;
mem[1*(ADDR_WIDTH)+67] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+68] =  32'b00110000000000010000000000000010;
mem[1*(ADDR_WIDTH)+69] =  32'b00110100100000010000000000000000;
mem[1*(ADDR_WIDTH)+70] =  32'b00110000000000010000000000001000;
mem[1*(ADDR_WIDTH)+71] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+72] =  32'b00110000000000010000000000000010;
mem[1*(ADDR_WIDTH)+73] =  32'b00110100100000010000000000000000;
mem[1*(ADDR_WIDTH)+74] =  32'b00110000000000010000000000001001;
mem[1*(ADDR_WIDTH)+75] =  32'b00001100001001000000000000000000;
mem[1*(ADDR_WIDTH)+76] =  32'b00110000000000010000000000001001;
mem[1*(ADDR_WIDTH)+77] =  32'b00110100100000010000000000000000;
mem[1*(ADDR_WIDTH)+78] =  32'b00110000000000010000000000000000;
mem[1*(ADDR_WIDTH)+79] =  32'b00110100000000010000000000010100;
mem[1*(ADDR_WIDTH)+80] =  32'b00110000000000010000000000001010;
mem[1*(ADDR_WIDTH)+81] =  32'b00110100000000010000000000010101;
mem[1*(ADDR_WIDTH)+82] =  32'b10000100000000000000000000000010;
mem[1*(ADDR_WIDTH)+83] =  32'b00001111101000010000000000000000;
mem[1*(ADDR_WIDTH)+84] =  32'b00110100000000010000000000011000;
mem[1*(ADDR_WIDTH)+85] =  32'b00101100000000010000000000011000;
mem[1*(ADDR_WIDTH)+86] =  32'b10110100000000010000000000000000;
mem[1*(ADDR_WIDTH)+87] =  32'b10101100000000000000000010000000;
mem[1*(ADDR_WIDTH)+88] =  32'b00000000000000000000000000000000;
mem[1*(ADDR_WIDTH)+89] =  32'b10101100000000000000000011000000;
mem[1*(ADDR_WIDTH)+90] =  32'b00000000000000000000000000000000;
mem[1*(ADDR_WIDTH)+91] =  32'b00000100000000000000000000000000;


mem[2*(ADDR_WIDTH)+0] =  32'b00000000000000000000000000000000;
mem[2*(ADDR_WIDTH)+1] =  32'b00111000000000000000000000110001;
mem[2*(ADDR_WIDTH)+2] =  32'b00101100000000010000000000000000;
mem[2*(ADDR_WIDTH)+3] =  32'b00001100001001000000000000000000;
mem[2*(ADDR_WIDTH)+4] =  32'b00110000000000010000000000000000;
mem[2*(ADDR_WIDTH)+5] =  32'b00001100001000100000000000000000;
mem[2*(ADDR_WIDTH)+6] =  32'b00001100100000110000000000000000;
mem[2*(ADDR_WIDTH)+7] =  32'b01011100011000100000000000001011;
mem[2*(ADDR_WIDTH)+8] =  32'b00110000000000010000000000000001;
mem[2*(ADDR_WIDTH)+9] =  32'b00001100001111010000000000000000;
mem[2*(ADDR_WIDTH)+10] =  32'b00111111111000000000000000000000;
mem[2*(ADDR_WIDTH)+11] =  32'b00101100000000010000000000000000;
mem[2*(ADDR_WIDTH)+12] =  32'b00001100001001000000000000000000;
mem[2*(ADDR_WIDTH)+13] =  32'b00110000000000010000000000000001;
mem[2*(ADDR_WIDTH)+14] =  32'b00001100001000100000000000000000;
mem[2*(ADDR_WIDTH)+15] =  32'b00001100100000110000000000000000;
mem[2*(ADDR_WIDTH)+16] =  32'b01011100011000100000000000010101;
mem[2*(ADDR_WIDTH)+17] =  32'b00110000000000010000000000000001;
mem[2*(ADDR_WIDTH)+18] =  32'b00001100001111010000000000000000;
mem[2*(ADDR_WIDTH)+19] =  32'b00111111111000000000000000000000;
mem[2*(ADDR_WIDTH)+20] =  32'b00111000000000000000000000110001;
mem[2*(ADDR_WIDTH)+21] =  32'b00101100000000010000000000000000;
mem[2*(ADDR_WIDTH)+22] =  32'b00001100001001000000000000000000;
mem[2*(ADDR_WIDTH)+23] =  32'b00001111110111101111111111111101;
mem[2*(ADDR_WIDTH)+24] =  32'b00110111110111110000000000000010;
mem[2*(ADDR_WIDTH)+25] =  32'b00101100000000010000000000000000;
mem[2*(ADDR_WIDTH)+26] =  32'b00110111110000010000000000000001;
mem[2*(ADDR_WIDTH)+27] =  32'b00110111110001000000000000000000;
mem[2*(ADDR_WIDTH)+28] =  32'b00101100000000010000000000000000;
mem[2*(ADDR_WIDTH)+29] =  32'b00001100001001010000000000000000;
mem[2*(ADDR_WIDTH)+30] =  32'b00110000000000010000000000000001;
mem[2*(ADDR_WIDTH)+31] =  32'b00001100001000100000000000000000;
mem[2*(ADDR_WIDTH)+32] =  32'b00001100101000110000000000000000;
mem[2*(ADDR_WIDTH)+33] =  32'b00010000011000100000100000000000;
mem[2*(ADDR_WIDTH)+34] =  32'b00110100000000010000000101011011;
mem[2*(ADDR_WIDTH)+35] =  32'b00101100000000010000000101011011;
mem[2*(ADDR_WIDTH)+36] =  32'b00110100000000010000000000000000;
mem[2*(ADDR_WIDTH)+37] =  32'b10000100000000000000000000000010;
mem[2*(ADDR_WIDTH)+38] =  32'b00101111110001000000000000000000;
mem[2*(ADDR_WIDTH)+39] =  32'b00101111110000010000000000000001;
mem[2*(ADDR_WIDTH)+40] =  32'b00110100000000010000000000000000;
mem[2*(ADDR_WIDTH)+41] =  32'b00101111110111110000000000000010;
mem[2*(ADDR_WIDTH)+42] =  32'b00001111110111100000000000000011;
mem[2*(ADDR_WIDTH)+43] =  32'b00001111101000010000000000000000;
mem[2*(ADDR_WIDTH)+44] =  32'b00001100001000100000000000000000;
mem[2*(ADDR_WIDTH)+45] =  32'b00001100100000110000000000000000;
mem[2*(ADDR_WIDTH)+46] =  32'b00011000011000100000100000000000;
mem[2*(ADDR_WIDTH)+47] =  32'b00001100001111010000000000000000;
mem[2*(ADDR_WIDTH)+48] =  32'b00111111111000000000000000000000;
mem[2*(ADDR_WIDTH)+49] =  32'b10101100000000000000000001000000;
mem[2*(ADDR_WIDTH)+50] =  32'b00000000000000000000000000000000;
mem[2*(ADDR_WIDTH)+51] =  32'b10110000000000010000000000000000;
mem[2*(ADDR_WIDTH)+52] =  32'b00110100000000010000000000000001;
mem[2*(ADDR_WIDTH)+53] =  32'b00101100000000010000000000000001;
mem[2*(ADDR_WIDTH)+54] =  32'b00110100000000010000000000000000;
mem[2*(ADDR_WIDTH)+55] =  32'b10000100000000000000000000000010;
mem[2*(ADDR_WIDTH)+56] =  32'b00001111101000010000000000000000;
mem[2*(ADDR_WIDTH)+57] =  32'b00110100000000010000000000000001;
mem[2*(ADDR_WIDTH)+58] =  32'b00101100000000010000000000000001;
mem[2*(ADDR_WIDTH)+59] =  32'b10110100000000010000000000000000;
mem[2*(ADDR_WIDTH)+60] =  32'b10101100000000000000000010000000;
mem[2*(ADDR_WIDTH)+61] =  32'b00000000000000000000000000000000;
mem[2*(ADDR_WIDTH)+62] =  32'b10101100000000000000000011000000;
mem[2*(ADDR_WIDTH)+63] =  32'b00000000000000000000000000000000;
mem[2*(ADDR_WIDTH)+64] =  32'b00000100000000000000000000000000;

mem[3*(ADDR_WIDTH)+0] =  32'b00000000000000000000000000000000;
mem[3*(ADDR_WIDTH)+1] =  32'b00111000000000000000000000111001;
mem[3*(ADDR_WIDTH)+2] =  32'b00101100000000010000000000000000;
mem[3*(ADDR_WIDTH)+3] =  32'b00001100001001000000000000000000;
mem[3*(ADDR_WIDTH)+4] =  32'b00110000000000010000000000000010;
mem[3*(ADDR_WIDTH)+5] =  32'b00001100001000100000000000000000;
mem[3*(ADDR_WIDTH)+6] =  32'b00001100100000110000000000000000;
mem[3*(ADDR_WIDTH)+7] =  32'b01110000011000100000000000001011;
mem[3*(ADDR_WIDTH)+8] =  32'b00110000000000010000000000000001;
mem[3*(ADDR_WIDTH)+9] =  32'b00001100001111010000000000000000;
mem[3*(ADDR_WIDTH)+10] =  32'b00111111111000000000000000000000;
mem[3*(ADDR_WIDTH)+11] =  32'b00001111110111101111111111111110;
mem[3*(ADDR_WIDTH)+12] =  32'b00110111110111110000000000000001;
mem[3*(ADDR_WIDTH)+13] =  32'b00101100000000010000000000000000;
mem[3*(ADDR_WIDTH)+14] =  32'b00110111110000010000000000000000;
mem[3*(ADDR_WIDTH)+15] =  32'b00101100000000010000000000000000;
mem[3*(ADDR_WIDTH)+16] =  32'b00001100001001000000000000000000;
mem[3*(ADDR_WIDTH)+17] =  32'b00110000000000010000000000000001;
mem[3*(ADDR_WIDTH)+18] =  32'b00001100001000100000000000000000;
mem[3*(ADDR_WIDTH)+19] =  32'b00001100100000110000000000000000;
mem[3*(ADDR_WIDTH)+20] =  32'b00010000011000100000100000000000;
mem[3*(ADDR_WIDTH)+21] =  32'b00110100000000010000000101011011;
mem[3*(ADDR_WIDTH)+22] =  32'b00101100000000010000000101011011;
mem[3*(ADDR_WIDTH)+23] =  32'b00110100000000010000000000000000;
mem[3*(ADDR_WIDTH)+24] =  32'b10000100000000000000000000000010;
mem[3*(ADDR_WIDTH)+25] =  32'b00101111110000010000000000000000;
mem[3*(ADDR_WIDTH)+26] =  32'b00110100000000010000000000000000;
mem[3*(ADDR_WIDTH)+27] =  32'b00101111110111110000000000000001;
mem[3*(ADDR_WIDTH)+28] =  32'b00001111110111100000000000000010;
mem[3*(ADDR_WIDTH)+29] =  32'b00001111101000010000000000000000;
mem[3*(ADDR_WIDTH)+30] =  32'b00001100001001000000000000000000;
mem[3*(ADDR_WIDTH)+31] =  32'b00001111110111101111111111111101;
mem[3*(ADDR_WIDTH)+32] =  32'b00110111110111110000000000000010;
mem[3*(ADDR_WIDTH)+33] =  32'b00101100000000010000000000000000;
mem[3*(ADDR_WIDTH)+34] =  32'b00110111110000010000000000000001;
mem[3*(ADDR_WIDTH)+35] =  32'b00110111110001000000000000000000;
mem[3*(ADDR_WIDTH)+36] =  32'b00101100000000010000000000000000;
mem[3*(ADDR_WIDTH)+37] =  32'b00001100001001010000000000000000;
mem[3*(ADDR_WIDTH)+38] =  32'b00110000000000010000000000000010;
mem[3*(ADDR_WIDTH)+39] =  32'b00001100001000100000000000000000;
mem[3*(ADDR_WIDTH)+40] =  32'b00001100101000110000000000000000;
mem[3*(ADDR_WIDTH)+41] =  32'b00010000011000100000100000000000;
mem[3*(ADDR_WIDTH)+42] =  32'b00110100000000010000000101011011;
mem[3*(ADDR_WIDTH)+43] =  32'b00101100000000010000000101011011;
mem[3*(ADDR_WIDTH)+44] =  32'b00110100000000010000000000000000;
mem[3*(ADDR_WIDTH)+45] =  32'b10000100000000000000000000000010;
mem[3*(ADDR_WIDTH)+46] =  32'b00101111110001000000000000000000;
mem[3*(ADDR_WIDTH)+47] =  32'b00101111110000010000000000000001;
mem[3*(ADDR_WIDTH)+48] =  32'b00110100000000010000000000000000;
mem[3*(ADDR_WIDTH)+49] =  32'b00101111110111110000000000000010;
mem[3*(ADDR_WIDTH)+50] =  32'b00001111110111100000000000000011;
mem[3*(ADDR_WIDTH)+51] =  32'b00001111101000010000000000000000;
mem[3*(ADDR_WIDTH)+52] =  32'b00001100001000100000000000000000;
mem[3*(ADDR_WIDTH)+53] =  32'b00001100100000110000000000000000;
mem[3*(ADDR_WIDTH)+54] =  32'b00001000011000100000100000000000;
mem[3*(ADDR_WIDTH)+55] =  32'b00001100001111010000000000000000;
mem[3*(ADDR_WIDTH)+56] =  32'b00111111111000000000000000000000;
mem[3*(ADDR_WIDTH)+57] =  32'b00110000000000010000000000000100;
mem[3*(ADDR_WIDTH)+58] =  32'b00110100000000010000000000000001;
mem[3*(ADDR_WIDTH)+59] =  32'b00101100000000010000000000000001;
mem[3*(ADDR_WIDTH)+60] =  32'b00110100000000010000000000000000;
mem[3*(ADDR_WIDTH)+61] =  32'b10000100000000000000000000000010;
mem[3*(ADDR_WIDTH)+62] =  32'b00001111101000010000000000000000;
mem[3*(ADDR_WIDTH)+63] =  32'b00110100000000010000000000000001;
mem[3*(ADDR_WIDTH)+64] =  32'b00101100000000010000000000000001;
mem[3*(ADDR_WIDTH)+65] =  32'b10110100000000010000000000000000;
mem[3*(ADDR_WIDTH)+66] =  32'b10101100000000000000000010000000;
mem[3*(ADDR_WIDTH)+67] =  32'b00000000000000000000000000000000;
mem[3*(ADDR_WIDTH)+68] =  32'b10101100000000000000000011000000;
mem[3*(ADDR_WIDTH)+69] =  32'b00000000000000000000000000000000;
mem[3*(ADDR_WIDTH)+70] =  32'b00000100000000000000000000000000;


mem[4*(ADDR_WIDTH)+0] =  32'b00000000000000000000000000000000;
mem[4*(ADDR_WIDTH)+1] =  32'b00111000000000000000000000011111;
mem[4*(ADDR_WIDTH)+2] =  32'b00110000000000010000000000000001;
mem[4*(ADDR_WIDTH)+3] =  32'b00110100000000010000000000000010;
mem[4*(ADDR_WIDTH)+4] =  32'b00110000000000010000000000000000;
mem[4*(ADDR_WIDTH)+5] =  32'b00110100000000010000000000000011;
mem[4*(ADDR_WIDTH)+6] =  32'b10000000000000000000000000000011;
mem[4*(ADDR_WIDTH)+7] =  32'b00101100000000010000000000000011;
mem[4*(ADDR_WIDTH)+8] =  32'b00001100001001000000000000000000;
mem[4*(ADDR_WIDTH)+9] =  32'b00101100000000010000000000000001;
mem[4*(ADDR_WIDTH)+10] =  32'b00001100001000100000000000000000;
mem[4*(ADDR_WIDTH)+11] =  32'b00001100100000110000000000000000;
mem[4*(ADDR_WIDTH)+12] =  32'b01110000011000100000000000011100;
mem[4*(ADDR_WIDTH)+13] =  32'b00101100000000010000000000000000;
mem[4*(ADDR_WIDTH)+14] =  32'b00001100001001000000000000000000;
mem[4*(ADDR_WIDTH)+15] =  32'b00101100000000010000000000000010;
mem[4*(ADDR_WIDTH)+16] =  32'b00001100001000100000000000000000;
mem[4*(ADDR_WIDTH)+17] =  32'b00001100100000110000000000000000;
mem[4*(ADDR_WIDTH)+18] =  32'b00011000011000100000100000000000;
mem[4*(ADDR_WIDTH)+19] =  32'b00110100000000010000000000000010;
mem[4*(ADDR_WIDTH)+20] =  32'b00101100000000010000000000000011;
mem[4*(ADDR_WIDTH)+21] =  32'b00001100001001000000000000000000;
mem[4*(ADDR_WIDTH)+22] =  32'b00110000000000010000000000000001;
mem[4*(ADDR_WIDTH)+23] =  32'b00001100001000100000000000000000;
mem[4*(ADDR_WIDTH)+24] =  32'b00001100100000110000000000000000;
mem[4*(ADDR_WIDTH)+25] =  32'b00001000011000100000100000000000;
mem[4*(ADDR_WIDTH)+26] =  32'b00110100000000010000000000000011;
mem[4*(ADDR_WIDTH)+27] =  32'b00111000000000000000000000000111;
mem[4*(ADDR_WIDTH)+28] =  32'b00101100000000010000000000000010;
mem[4*(ADDR_WIDTH)+29] =  32'b00001100001111010000000000000000;
mem[4*(ADDR_WIDTH)+30] =  32'b00111111111000000000000000000000;
mem[4*(ADDR_WIDTH)+31] =  32'b10101100000000000000000001000000;
mem[4*(ADDR_WIDTH)+32] =  32'b00000000000000000000000000000000;
mem[4*(ADDR_WIDTH)+33] =  32'b10110000000000010000000000000000;
mem[4*(ADDR_WIDTH)+34] =  32'b00110100000000010000000000000101;
mem[4*(ADDR_WIDTH)+35] =  32'b10101100000000000000000001000000;
mem[4*(ADDR_WIDTH)+36] =  32'b00000000000000000000000000000000;
mem[4*(ADDR_WIDTH)+37] =  32'b10110000000000010000000000000000;
mem[4*(ADDR_WIDTH)+38] =  32'b00110100000000010000000000000110;
mem[4*(ADDR_WIDTH)+39] =  32'b00101100000000010000000000000101;
mem[4*(ADDR_WIDTH)+40] =  32'b00110100000000010000000000000000;
mem[4*(ADDR_WIDTH)+41] =  32'b00101100000000010000000000000110;
mem[4*(ADDR_WIDTH)+42] =  32'b00110100000000010000000000000001;
mem[4*(ADDR_WIDTH)+43] =  32'b10000100000000000000000000000010;
mem[4*(ADDR_WIDTH)+44] =  32'b00001111101000010000000000000000;
mem[4*(ADDR_WIDTH)+45] =  32'b00110100000000010000000000000100;
mem[4*(ADDR_WIDTH)+46] =  32'b00101100000000010000000000000100;
mem[4*(ADDR_WIDTH)+47] =  32'b10110100000000010000000000000000;
mem[4*(ADDR_WIDTH)+48] =  32'b10101100000000000000000010000000;
mem[4*(ADDR_WIDTH)+49] =  32'b00000000000000000000000000000000;
mem[4*(ADDR_WIDTH)+50] =  32'b10101100000000000000000011000000;
mem[4*(ADDR_WIDTH)+51] =  32'b00000000000000000000000000000000;
mem[4*(ADDR_WIDTH)+52] =  32'b00000100000000000000000000000000;*/


	end
	
	always @ (posedge clock)
		begin
			if( writeInstr )
				mem[(ADDR_WIDTH)*WritepId + HDAddress] <= instrIn;
		end
	always @( posedge autoclock )
		begin
			InstructionOut <= mem[(ADDR_WIDTH)*region + address];
		end
endmodule
	