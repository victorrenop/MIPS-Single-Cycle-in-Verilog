module InstructionMemory (adress, InstructionOut, clock);

	input [9:0] adress;
	input clock;
	output [31:0] InstructionOut;
	reg [31:0] mem [55:0];
	integer flag = 0;
	
	always @ (posedge clock)
		begin
			if (flag == 0)
			begin
				
				/*
				//Fibonacci
				mem[0] = 32'b00000000000000000000000000000000; // nop
				mem[1] = 32'b00110000000001100000000000000000; // r[6] = Im(0)
				mem[2] = 32'b00110000000001110000000000000001; // r[7] = Im(1)
				mem[3] = 32'b01111100000000010000000000000000; // in reg[1]
				mem[4] = 32'b00010100001000010000000000000001; // r[1] = r[1] - Im(1)
				mem[5] = 32'b00110000000000100000000000000001; // r[2] = Im(1)
				mem[6] = 32'b00110000000000110000000000000000; // r[3] = Im(0)
				mem[7] = 32'b01101100011000010000000000010011; // r[3] > r[1], PC = 19
				mem[8] = 32'b01101100011000100000000000001100; // r[3] > r[2], PC = 12
				mem[9] = 32'b00001000011000000010100000000000; // r[5] = r[3] + r[0]
				mem[10] = 32'b00110100000001010000000000000001; // MEM[r[0] + Im(1)] = r[5]
				mem[11] = 32'b00111000000000000000000000010000; // PC = 16
				mem[12] = 32'b00001000110001110010100000000000; // r[5] = r[6] + r[7]
				mem[13] = 32'b00001000111000000011000000000000; // r[6] = r[7] + r[0]
				mem[14] = 32'b00001000101000000011100000000000; // r[7] = r[5] + r[0]
				mem[15] = 32'b00110100000001010000000000000001; // MEM[r[0] + Im(1)] = r[5]
				mem[16] = 32'b10000000000000000000000000000001; // out reg[1]
				mem[17] = 32'b00001100011000110000000000000001; // r[3] = r[3] + Im(1)
				mem[18] = 32'b00111000000000000000000000000111; // PC = 7
				mem[19] = 32'b00101100000010110000000000000001; // r[11] = MEM[r[0] + Im(1)]	
				mem[20] = 32'b00010101011010110000000000000010; // r[11] = r[11] - Im(1)
				mem[21] = 32'b00110100000010110000000000000010; // MEM[r[0] + Im(2)] = r[11]
				mem[22] = 32'b10000000000000000000000000000010; // out reg[2]
				
				
				
				//Insertion Sort
				mem[0] = 32'b00000000000000000000000000000000; // nop
				mem[1] = 32'b01111100000000010000000000000000; // in reg[1]
				mem[2] = 32'b00110000000000110000000000000001; // r[3] = Im(1)
				mem[3] = 32'b00110000000001000000000000001100; // r[4] = Im(12)
				mem[4] = 32'b00110000000001010000000000001111; // r[5] = Im(15)
				mem[5] = 32'b00110000000001100000000000000110; // r[6] = Im(6)
				mem[6] = 32'b00110000000001110000000000001010; // r[7] = Im(10)
				mem[7] = 32'b00110000000010000000000000000001; // r[8] = Im(1)
				mem[8] = 32'b00110000000010010000000000000000; // r[9] = Im(0)
				mem[9] = 32'b00110000000000100000000000100101; // r[2] = Im(37)
				mem[10] = 32'b00110100000000100000000000000001; // MEM[r[0] + Im(1)] = r[2]
				mem[11] = 32'b00110100000000110000000000000010; // MEM[r[0] + Im(2)] = r[3]
				mem[12] = 32'b00110100000001000000000000000011; // MEM[r[0] + Im(3)] = r[4]
				mem[13] = 32'b00110100000001010000000000000100; // MEM[r[0] + Im(4)] = r[5]
				mem[14] = 32'b00110100000001100000000000000101; // MEM[r[0] + Im(5)] = r[6]
				mem[15] = 32'b00110100000001110000000000000110; // MEM[r[0] + Im(6)] = r[7]
				mem[16] = 32'b01101101000000010000000000011101; // r[8] > r[1], PC = 29
				mem[17] = 32'b00010101000010010000000000000001; // r[9] = r[8] - Im(1)
				mem[18] = 32'b00101101000010100000000000000000; // r[10] = MEM[r[8] + Im(0)]
				
				mem[19] = 32'b01111001001000000000000000011010; // r[9] < r[0], PC = 26
				
				mem[20] = 32'b00101101001011000000000000000000; // r[12] = MEM[r[9] + Im(0)]
				mem[21] = 32'b01101101010011000000000000011010; // r[10] > r[12], PC = 26
				mem[22] = 32'b00101101001010110000000000000000; // r[11] = MEM[r[9] + Im(0)]
				mem[23] = 32'b00110101001010110000000000000001; // MEM[r[9] + Im(1)] = r[11]
				mem[24] = 32'b00010101001010010000000000000001; // r[9] = r[9] - Im(1)
				mem[25] = 32'b00111000000000000000000000010011; // PC = 19
				
				mem[26] = 32'b00110101001010100000000000000001; // MEM[r[9] + Im(1)] = r[10]
				mem[27] = 32'b00001101000010000000000000000001; // r[8] = r[8] + Im(1)
				mem[28] = 32'b00111000000000000000000000010000; // PC = 16
				mem[29] = 32'b10000000000000000000000000000001; // out reg[1]
				mem[30] = 32'b10000000000000000000000000000010; // out reg[2]
				mem[31] = 32'b10000000000000000000000000000011; // out reg[3]
				mem[32] = 32'b10000000000000000000000000000100; // out reg[4]
				mem[33] = 32'b10000000000000000000000000000101; // out reg[5]
				mem[34] = 32'b10000000000000000000000000000110; // out reg[6]
				mem[35] = 32'b10000000000000000000000000000111; // out reg[7]
				*/
				
				
				//Todas as instrcoes
				mem[0] = 32'b00000000000000000000000000000000; // nop
				mem[1] = 32'b01111100000000010000000000000000; // in reg[1]
				mem[2] = 32'b00110000000000100000000000000111; // r[2] = Im(7)
				mem[3] = 32'b00001000001000100001100000000000; // r[3] = r[1] + r[2]
				mem[4] = 32'b00001100001001000000000000001101; // r[4] = r[1] + Im(13)
				mem[5] = 32'b00010000001000100010100000000000; // r[5] = r[1] - r[2]
				mem[6] = 32'b00010100100001100000000000000111; // r[6] = r[4] - Im(7)
				mem[7] = 32'b00011000001000100100000000000000; // r[8] = r[1] * r[2]
				mem[8] = 32'b00011101000001000100100000000000; // r[9] = r[8] / r[4]
				mem[9] = 32'b00100000001000100011100000000000; // r[7] = r[1] < r[2]
				mem[10] = 32'b00100100100010110000000001000000; // r[11] = r[4] >> 1
				mem[11] = 32'b00101001000011000000000001000000; // r[12] = r[8] << 1
				mem[12] = 32'b00110100000010000000000000000001; // MEM[r[0] + Im(1)] = r[8]
				mem[13] = 32'b00101100000010110000000000000001; // r[11] = MEM[r[0] + Im(1)]
				mem[14] = 32'b10000000000000000000000000000001; // out reg[1]
				mem[15] = 32'b00110100000000110000000000000010; // MEM[r[0] + Im(2)] = r[3]
				mem[16] = 32'b10000000000000000000000000000010; // out reg[2]
				mem[17] = 32'b00111000000000000000000000011110; // PC = 30
				mem[30] = 32'b01000000001000100110100000000000; // r[13] = r[1] ^ r[2]
				mem[31] = 32'b01000100001000100111000000000000; // r[14] = r[1] && r[2]
				mem[32] = 32'b01001000001000110111100000000000; // r[15] = r[1] || r[3]
				mem[33] = 32'b01001100001100000000000000000000; // r[16] = ~r[1]
				mem[34] = 32'b01010000001100010000000000001101; // r[17] = r[1] ^ Im(13)
				mem[35] = 32'b01010100001100100000000000001101; // r[18] = r[1] && Im(13)
				mem[36] = 32'b01011000001100110000000000001101; // r[19] = r[1] || Im(13)
				mem[37] = 32'b01111100000101000000000000000000; // in reg[20]
				mem[38] = 32'b01011100001101000000000000101000; // r[1] == r[20], PC = 40
				mem[40] = 32'b00000000000000000000000000000000; // nop
				mem[41] = 32'b01101000001000000000000000110001;// r[1] != r[0], PC = 49
				mem[44] = 32'b01110000001000100000000000101111; // r[1] < r[2], PC = 47
				mem[47] = 32'b01110100001000000000000000110011; // r[1] > r[0], PC = 51
				mem[49] = 32'b01101100010000010000000000101100; // r[2] > r[1], PC = 44
				mem[51] = 32'b01111000101000000000000000110111; // r[5] < r[0], PC = 55
				mem[55] = 32'b10000000000000000000000000000001; // out reg[1]	
				
				
				flag <= 1;
			end
		end	
		assign InstructionOut = mem[adress];
endmodule
	